ab	ab
abba	abba
abbas	abbas
abbey	abbey
abc	abc
abort	abortion
aborter	abortions
about	about
abraham	abraham
absint	absinthe
absolut	absolute
absoluta	absolute
absolution	absolution
absorberas	(gets) absorbed
abstrakta	abstract
abu	abu
ac	ac
academy	academy
acceptera	accept
accepterad	accepted
accepterade	accepted
accepterar	accept
accepterat	accepted
acdc	ac/dc
action	action
ad	ad
adam	adam
adams	adams
adeln	nobility
adhd	adhd
adjektiv	adjective
administration	administration
administrationen	administration
administrativ	administrative
administrativa	administrative
administrativt	administratively
adolf	adolf
adolfs	adolf
adrian	adrian
advokat	lawyer
af	of (old swedish)
affärer	business
afghanistan	afghanistan
africa	africa
afrika	africa
afrikaner	africans
afrikansk	african
afrikanska	african
afrikas	africa
afrodite	afrodite
aftonbladet	aftonbladet
age	age
agent	agent
agera	act
agerande	behavior
aggressiv	aggressive
agnes	agnes
agnetha	agnetha
agnosticism	agnosticism
agnostiker	agnostic
ahmed	ahmed
aids	aids
aik	aik
airlines	airlines
airport	airport
ajax	ajax
akademi	academy
akademien	academy
akademiens	academy
akademisk	academic
akademiska	academic
akc	akc
akon	akon
akondroplasi	achondroplasia
aktiebolag	companies
aktier	stock
aktiv	active
aktiva	active
aktivitet	activity
aktiviteten	activity
aktiviteter	activities
aktivt	active
aktuell	current
aktuella	current
aktuellt	current
aktörer	actors
akut	acute
al	alder
alan	alan
alaska	alaska
albaner	albanians
albanien	albania
albanska	albanian
albert	albert
album	album
albumen	album
albumet	album
albumets	album
alces	alces
aldrig	never
ale	ale
alex	alex
alexander	alexander
alexanders	alexanders
alexandra	alexandra
alexandria	alexandria
alf	alf
alfa	alpha
alfabet	alphabet
alfabetet	alphabet
alfabetisk	alphabetical
alfred	alfred
alger	algaes
algeriet	algeria
ali	ali
alice	alice
alkohol	alcohol
alkoholer	alcohols
alla	all
allan	allan
alldeles	right
allen	allen
allians	alliance
alliansen	alliance
allierad	ally
allierade	allied
allierades	allied
allmän	general
allmänhet	public
allmänheten	public
allmänna	general
allmänt	generally
allra	very
alls	all
allsvenskan	allsvenskan
allt	all
alltför	all too
alltid	always
allting	everything
alltjämt	still
alltmer	increasingly
alltsedan	since
alltså	so
allvar	earnest
allvarlig	serious
allvarliga	serious
allvarligt	serious
alperna	alps
alqaida	al-qaida
alternativ	alternative
alternativa	alternative
alternativt	alternatively
aluminium	aluminum
am	am
amazonas	the amazon rainforest
ambassad	embassy
ambitioner	ambitions
america	america
american	american
amerika	america
amerikanen	american
amerikaner	americans
amerikanerna	americans
amerikansk	american
amerikanska	us
amerikanske	american
amerikanskt	american
amerikas	america
amfetamin	amphetamine
aminosyra	amino acid
aminosyror	amino acids
ammoniak	ammonia
amsterdam	amsterdam
amy	amy
ana	feel
analsex	anal sex
analys	analysis
analytisk	analytical
analytiska	analytical
anarkism	anarchism
anarkismen	anarchism
anarkister	anarchists
anarkistiska	anarchistic
anatolien	anatolia
anatomi	anatomy
anc	anc
anda	spirit
andas	breath
ande	spirit
andel	share
andelen	share
anden	spirit
anderna	andes
anders	anders
andersson	andersson
anderssons	andersson
andlig	spiritual
andliga	spiritual
andra	other
andras	others
andre	second
andreas	andreas
andres	andres
andrew	andrew
andré	andre
andy	andy
anfall	attack
anfalla	attack
anfallet	attack
anfield	anfield
anföll	attacked
ange	set
angeles	angeles
angelina	angelina
angels	angels
anger	indicates
anges	out
anglosaxiska	anglo-saxon
angola	angola
angrepp	attack
angränsande	adjacent
angående	concerning
anhängare	supporters
anhöriga	kin
animerade	animated
anka	duck
anklagade	accused
anklagades	accused
anklagats	accused
anklagelser	accusations
anknytning	connection
ankomst	arrival
anlades	were built
anledning	reason
anledningar	reasons
anledningarna	reasons
anledningen	reason
anläggningar	plants
anlände	arrived
anländer	arrives
anna	anna
annan	other
annars	else
annat	other
anne	anne
annekterade	annexed
annika	amy
annorlunda	different
anor	ancestry
anordnas	provided
anorektiker	anorectics
anorexia	anorexia
another	another
anpassa	adapt
anpassade	custom
anpassat	adapted
anpassning	adaption
anser	view
anses	considered
ansetts	considered
ansikte	face
ansiktet	face
ansluta	connect
ansluter	connects
anslutna	connected
anslutning	connection
anslöt	joined
anspråk	claim
ansträngningar	effort
anställd	employed
anställda	employees
ansvar	responsibility
ansvarar	responsible
ansvaret	responsibility
ansvarig	responsible
ansvariga	responsible
ansåg	felt
ansågs	was
ansökte	applied
anta	adopting
antagit	adopted
antagits	adoption
antagligen	probably
antal	number of
antalet	number
antar	suppose
antarktis	antarctica
antarktiska	antarctic
antas	adoption
anteckningar	notes
anthony	anthony
antika	old
antiken	the ancient world
antikens	ancient
antingen	either
antisemitiska	antisemitic
antisemitism	antisemitism
antisemitismen	antisemitism
antog	adopted
antogs	adopted
antoinette	antoinette
antonio	antonio
antropogen	anthropogenic
antyder	indicates
anus	anus
använda	use
användande	using
användandet	use
användare	user
användaren	user
användas	used
användbar	useful
användbara	useful
använder	using
användes	used
användning	use
användningen	use
användningsområden	applications
används	used
använt	used
använts	used
apartheid	apartheid
apollo	apollo
april	april
ar	is
arab	arab
arabemiraten	uae
araber	arab
araberna	arabs
arabisk	arab
arabiska	arabic
arabvärlden	arab
arbeta	work
arbetade	worked
arbetar	working
arbetare	workers
arbetarklassen	working
arbetat	worked
arbete	work
arbeten	works
arbetet	the work
arbetsgivare	employer
arbetsgivaren	employer
arbetskraft	workforce
arbetslöshet	unemployment
arbetslösheten	unemployment
arbetsplats	workplace
area	area
arean	area
arena	arena
arenan	arena
arg	angry
argentina	argentina
argument	argument
aristokratin	nobility
aristoteles	aristotle
arkeologiska	archaeological
arkitekt	architect
arkitekten	architect
arkitekter	architects
arkitektur	architecture
arkitekturen	architecture
arkiv	archive
arlanda	arlanda
arm	arm
armar	arms
armenien	armenian
armeniska	armenian
army	army
armé	army
arméer	armies
arméerna	armies
armén	army
arméns	army
arnold	arnold
arrangemang	arrangement
arrangeras	arranged
arresterades	was arrested
arsenal	arsenal
art	species
arten	species
arter	species
arterna	species
arternas	species
arthur	arthur
artikel	article
artikeln	the article
artiklar	items
artist	artist
artisten	artist
artister	artists
artisterna	performers
arton	eighteen
arvet	the inheritance
arvid	arvid
asiatiska	asian
asien	asia
aspekt	aspect
aspekter	aspects
aspergers	aspergers
assistent	assistant
assisterande	assistant
assyriska	assyrian
asterix	asterix
asteroidbältet	the asteroid belt
asteroider	asteroids
aston	aston
astrid	astrid
astronomer	astronomers
astronomi	astronomy
astronomin	astronomy
astronomiska	astronomical
ateism	atheism
ateist	atheist
ateister	atheists
aten	general
atlanta	atlanta
atlanten	atlantic
atlas	atlas
atmosfär	atmosphere
atmosfären	atmosphere
atom	atom
atombomben	atomic bomb
atombomberna	atomic bomb
atomer	atoms
atomkärnor	nuclei
att	to
attacken	attack
attacker	attacks
attackerna	attacks
august	august
augusti	august
auktoritet	authority
auktoritära	authoritarian
auschwitz	auschwitz
austin	austin
australia	australia
australian	australian
australien	australia
australiens	australia
australiska	australian
autism	autism
automatiskt	automatic
autonom	autonomous
autonoma	autonomous
autonomi	autonomy
av	of
avalanche	avalanche
avancerad	advanced
avancerade	advanced
avbrott	break
avbryta	cancel
avbröts	canceled
avel	breeding
avfall	waste
avgick	resigned
avgå	resign
avgör	decides
avgöra	determine
avgörande	settling
avgörs	determined
avhandling	thesis
avkomma	offspring
avled	died
avlidit	dies
avlidna	deceased
avlägsna	remove
avrättades	executed
avrättning	execution
avrättningar	executions
avrättningen	execution
avsaknad	lack
avsaknaden	lack
avsattes	deposited
avsedd	intended
avsedda	intended
avseende	respect
avseenden	regard
avser	refers
avses	referred
avsett	intended
avsevärt	considerably
avsikt	intention
avsikten	intent
avskaffa	abolish
avskaffade	abolished
avskaffades	abolished
avskaffande	abolition
avskaffandet	abolition
avsluta	end
avslutade	finished
avslutades	completed
avslutas	ends
avslutat	finished
avslöjade	revealed
avsnitt	episode
avsnitten	the episodes
avsnittet	section
avstå	refrain
avstånd	distance
avståndet	distance
avsätta	unseat
avsåg	related
avtal	agreement
avtalet	agreement
avtar	decreases
avvikande	different
avvikelser	deviations
avvisade	rejected
avvisar	reject
awards	awards
axel	axel
axelmakterna	axis
axl	axl
azerbajdzjan	azerbaijan
azidgrupp	azide group
b	b
babylon	babylon
bad	swimming
bagge	ram
bahamas	bahamas
baháulláh	bahullah
baháí	bahá'í
baker	baker
bakgrund	background
bakom	behind
bakterier	bacteria
bakåt	backwards
balans	balance
balansen	balance
balkan	the balkans
balkanhalvön	balkan peninsula
baltikum	baltics
baltimore	baltimore
baltiska	baltic
bana	course
banan	banana
banbrytande	groundbreaking
band	band
banden	bander
bandet	band
bandets	band
bandmedlemmar	band members
bandmedlemmarna	band members
bank	bank
banker	banks
banor	paths
baptism	baptist
bar	bar
bara	only
barack	barracks
barbro	barbro
barcelona	barcelona
barcelonas	barcelona
barndom	childhood
barnen	children
barnens	children
barnet	child
barnets	child
barney	barney
barns	child
baron	baron
barrett	barrett
barry	barry
bars	bar
bart	offense
bas	base
basen	base
baser	bases
baserad	based
baserade	based
baserar	base
baseras	based
baserat	based
basis	basis
basist	bassist
basisten	bassist
basket	basketball
batman	batman
bay	bay
bayern	bayern
bbc	bbc
be	ask
beatles	beatles
bebott	inhabited
bebyggelse	buildings
bebyggelsen	buildings
beck	pitch
beckham	beckham
bedrev	conducted
bedriva	carry
bedriver	manage
bedrivs	conducted
bedöma	judge; decide
bedöms	expected
beethoven	beethoven
befann	found
befinna	be
befinner	is
befintliga	existing
befogenhet	authority
befogenheter	powers
befolkade	populated
befolkning	population
befolkningen	population
befolkningens	population
befolkningstillväxt	population growth
befolkningstillväxten	population growth
befolkningstäthet	population density
befolkningstätheten	population density
befolkningsutveckling	demographics
befruktning	fertilization
befäl	command
befälet	command
befälhavare	commander
begav	went
begick	committed
begravd	buried
begravdes	buried
begravning	funeral
begrepp	concept
begreppen	the concepts
begreppet	the concept
begränsa	limit
begränsad	limited
begränsade	limited
begränsar	limit
begränsas	restricted
begränsat	restricted
begränsningar	limitations
begär	asks
begäran	request
begärde	called
begå	commit
begår	commits
begått	committed
behandla	treat
behandlade	treated
behandlades	treated
behandlar	treat
behandlas	treated
behandling	treatment
behandlingar	treatments
behandlingen	treatment
behov	needs
behovet	need
behålla	retain
behåller	retain
behöll	kept
behöva	need
behövde	needed
behövdes	needed
behöver	requires
behövs	required
bekant	known
bekostnad	expense
bekräftade	confirmed
bekräftades	confirmed
bekräftar	confirms
bekräftat	confirmed
bekämpa	prevent
belagt	coated
belgien	belgium
belgiens	belgium
belgiska	belgian
belgrad	belgrade
bell	bell
bella	bella
belopp	amount
belägen	located
beläget	located
belägg	evidence
belägna	located
belönades	awarded
bemärkelse	sense
ben	bone
benen	legs
benfica	benfica
bengt	bengt
bengtsson	bengtsson
benny	benny
bensin	gasoline
benämnas	named
benämning	name
benämningar	terms
benämningen	designation
benämns	designated
beordrade	ordered
ber	asks
beredd	prepared
berg	mountain
bergarter	rocks
bergen	mountain
berger	berger
berget	mount
bergman	bergman
bergmans	bergman
bergqvist	bergqvist
bergskedjan	mountain range
bergskedjor	mountain ranges
berlin	berlin
berlinmuren	berlin
berlins	berlin
bernadotte	bernadotte
bernhard	bernhard
bero	depend
berodde	was
beroende	dependent
beroendeframkallande	addictive
beror	depend
bertil	bertil
beräkna	calculate
beräknades	calculated
beräknar	computes
beräknas	calculated
beräkningar	calculations
berätta	tell
berättade	told
berättar	says
berättas	told
berättat	told
berättelse	story
berättelsen	story
berättelser	stories
berättelserna	stories
berömd	famous
berömda	famous
berömt	famous
berör	affecting
besegra	defeat
besegrade	defeated
besegrades	defeated
besegrat	defeated
besittning	possess
besittningar	holdings
beskrev	described
beskrevs	described
beskriva	describe
beskrivas	described
beskriver	describes
beskrivit	described
beskrivits	described
beskrivning	description
beskrivningar	descriptions
beskrivningen	description
beskrivs	described
beskydd	protection
beskyddare	patron
beslut	decision
beslutade	decided
beslutar	decides
beslutat	decided
besluten	decisions
beslutet	decision
besläktade	related
besläktat	related
beslöt	decided
besserwisser	wiseacre
best	best
bestod	was
bestämd	determined
bestämde	decided
bestämdes	determined
bestämma	determine
bestämmelser	regulations
bestämmer	decide
bestäms	determined
bestämt	certainly
bestå	consists
bestående	comprising
beståndsdelar	ingredients
består	consists
besättningen	crew
besök	visit
besöka	visit
besökare	visitors
besöker	visit
besökt	visit
besökte	visited
bet	bit
beta	beta
betala	pay
betalade	payed
betalar	pay
betalt	charge
beteckna	designate
betecknar	represents
betecknas	designated
beteckning	designation
beteckningen	designation
beteende	behavior
beteenden	behavior
betonade	emphasized
betonar	stress
betoning	stress
betrakta	regard
betraktade	observed
betraktades	considered
betraktar	regard
betraktas	considered
betraktats	considered
betyda	mean
betydande	important
betydde	meant
betydelse	meaning
betydelsefull	important
betydelsefulla	significant
betydelsen	meaning
betydelser	meanings
betyder	mean
betydligt	considerably
betyg	grade
bevara	preserve
bevarad	preserved
bevarade	preserved
bevaras	preserved
bevarat	preserved
bevarats	preserved
bevis	evidence
bevisa	prove
beväpnade	armed
beyoncé	beyoncé
bibel	bible
bibeln	bible
bibelns	bible
bibliografi	bibliography
bibliotek	library
bibliska	biblican
bidra	contribute
bidrag	contribution
bidragande	contributors
bidragen	the contributions
bidraget	grant
bidragit	contributed
bidrar	help
bidrog	contributed
big	big
bil	car
bilar	cars
bilbo	bilbo
bild	picture
bilda	form
bildade	formed
bildades	formed
bildande	formation
bildandet	formation
bildar	form
bildas	formed
bildat	formed
bildats	formed
bilden	image
bilder	pictures
bilderna	the pictures
bildning	formation
bildt	bildt
bilen	car
billboardlistan	bilboardlist
billiga	cheap
billy	billy
bilmärke	car make
binda	bind
bindande	binding
binder	bind
binds	bound
bioetik	bioethics
biogeografi	biogeography
biografen	the cinema
biografer	cinemas
biografi	biography
biologi	biology
biologisk	biological
biologiska	biological
bipolär	bipolar
bipolära	bipolar
birger	birger
birgitta	birgitta
birk	birk
birmingham	birmingham
biskop	bishop
biskopen	bishop
bistånd	aid
bit	bit
bitar	pieces
biträdande	assistant
bitter	bitter
bjöd	commanded
björn	björn
bl	inter
bla	blah
black	black
blad	leaf
blanc	blanc
bland	inter
blanda	mix
blandad	mixed
blandade	mixed
blandas	mixed
blandat	mixed
blandning	mixture
blekinge	blekinge
blev	became
bli	become
blind	blind
blir	gets
blivande	future
blivit	been
block	block
blod	blood
blodet	blood
blodiga	bloody
blodkroppar	corpuscle
blodtryck	blood pressure
blodtrycket	blood pressure
blogg	blog
bloggar	blogs
blommor	flowers
blomstrade	flourished
blott	only
blue	blue
blues	blues
bly	lead
bläckpenna	pen
blå	blue
blåser	blowing
blått	blue
blåvitt	blåvitt
bmi	bmi
bnp	gdp
bob	bob
bobby	bobby
bodde	lived
boende	resident
bojkott	boycott
bok	book
boken	the book
bokförlaget	publishing
bokstav	letter
bokstaven	the letter
bokstäver	letters
bokstäverna	letters
bolag	company
bolaget	company
bolagets	company
bolivia	bolivia
bolivianska	bolivian
bolivias	bolivia
bollen	ball
bolsjevikerna	the bolsheviks
bolt	bolt
bomb	bomb
bomben	bomb
bomber	bombs
bomull	cotton
bon	bon
bonaparte	bonaparte
bond	bond
bonde	farmer
bonniers	bonniers
book	book
bor	live
bord	table
borde	should
bordet	table
borg	castle
borgen	bail
borgerliga	civil
borgmästare	mayor
boris	boris
born	born
borrelia	borrelia
bort	away
borta	away
bortgång	death
bortom	beyond
bortsett	except
bosatt	resident
bosatta	residents
bosatte	settled
bosnien	bosnia
bosnienhercegovina	bosnia-hercegovina
bostad	residence
bostadsområden	residential
boston	boston
bostäder	housing
bosättare	settlers
bosättningar	settlements
bott	stayed
botten	bottom
bowie	bowie
boxning	boxing
boy	boy
bra	good
brad	brad
brand	fire
branden	fire
brandenburg	brandenburg
brasilianska	brasilian
brasilien	brazil
brasiliens	brazil
breaking	breaking
bred	wide
breda	broad
bredare	wider
breddgraden	parallel
bredvid	beside
brev	letter
brevet	the letter
brian	brian
bridge	bridge
brinnande	burning
brinner	on fire
brist	lack
bristande	lack
bristen	lack
brister	inabilities
brita	brita
britannica	britannica
british	british
britney	britney
britter	british
britterna	british
brittisk	british
brittiska	british
brittiske	british
brittiskt	british
bro	bridge
broar	bridges
broder	brother
brodern	brother
bron	bridge
brons	bronze
bronsåldern	bronze age
bronx	bronx
brooke	brooke
brooklyn	brooklyn
bror	brother
brother	brother
brott	crime
brottet	offense
brottslighet	crime
brottslingar	criminals
brown	brown
bruce	bruce
bruk	use
brukade	used
brukar	usually
bruket	the use
brushane	ruff
brutit	broken
bruttonationalprodukt	gdp
bryssel	brussels
bryta	break
bryter	breaking
bryts	broken
bränder	fires
brändes	burnt
brännvin	schnaps
bränsle	fuel
bränslen	fuel
bråk	brawl; fight
bröd	bread
bröder	brothers
bröderna	brothers
bröllop	wedding
bröllopet	wedding
bröstet	breast
bröt	broke
bröts	broken
bud	bid
budapest	budapest
buddha	buddha
buddhas	buddha
buddhism	buddhism
buddhismen	buddhism
buddhister	buddhist
buddhistiska	buddhist
buddy	buddy
budet	bid
budget	budget
budgeten	budget
budskap	message
budskapet	message
bulgarien	bulgaria
bulgariens	bulgaria
bulgariska	bulgarian
bundna	bound
bunny	bunny
burj	burj
burma	burma
burr	burr
burton	burton
burundi	burundi
bush	bush
bushadministrationen	bush administration
bushs	bush
buss	bus
bussar	bus
butiker	shops
by	village
byar	villages
bygga	build
byggandet	construction
byggas	prevented
byggd	built
byggda	built
byggde	built
byggdes	built
bygger	based
bygget	construction
byggnad	building
byggnaden	the building
byggnader	buildings
byggnaderna	buildings
byggnadsverk	building
byggs	built
byggt	built
byggts	built
byn	village
byrå	bureau
bysantinska	byzantine
byta	change
byte	change
byten	byte
byter	change
bytet	change
byts	changed
bytt	changed
bytte	changed
byttes	changed
byxor	pants
bägge	both
bär	carrying
bära	carry
bärande	carrying
bäst	best
bästa	top
bäste	best
bättre	better
båda	both
både	both
bål	prom
båt	boat
båtar	boats
båten	the boat
böcker	books
böckerna	books
böhmen	bohemia
bön	prayer
bönder	farmers
bönderna	farmers
bönor	beans
bönorna	beans
bör	should
bördiga	fertile
börja	start
började	started
början	beginning
börjar	begins
börjat	began
börje	borje
ca	cirka
caesar	caesar
caesars	caesar
café	coffeehouse
california	california
calle	calle
cambridge	cambridge
camp	camp
campus	campus
can	can
canada	canada
canadian	canadian
canaria	canaria
cancer	cancer
cannabis	cannabis
cant	cant
capita	head
capitol	capitol
carl	carl
carlo	carlo
carlos	carlos
carlsson	carlsson
carola	carola
carolina	carolina
carter	carter
cash	cash
casino	casino
castro	castro
cd	cd
cecilia	cecilia
cell	cell
cellen	cell
cellens	cell
celler	cells
cellerna	cells
census	census
center	center
centra	centers
central	central
centrala	central
centralamerika	central america
centralasien	central asia
centralbanken	central bank
centraleuropa	central
centralort	seat
centralorter	regional centers
centralstation	central
centralt	central
centre	center
centrum	center
champagne	champagne
chandler	chandler
channel	channel
chans	chance
chansen	chance
chaplin	chaplin
charles	charles
charlie	charlie
charlotte	charlotte
chefen	head
chelsea	chelsea
chi	chi
chicago	chicago
chile	chile
chiles	chile
chili	chili
choice	choice
choklad	chocolate
chokladen	chocolate
chris	chris
christer	christer
christian	christian
christina	christina
chrusjtjov	chrusjtjov
church	church
churchill	churchill
cia	cia
cirka	about
cirkel	circular
citat	quote
city	city
civil	civil
civila	civil
civilbefolkningen	civilians
civilisationen	civilization
civilisationer	civilizations
claes	claes
claude	claude
cliff	cliff
clinton	clinton
club	club
cobain	cobain
cocacola	coca-cola
cohen	cohen
coldplay	coldplay
colin	colin
colombia	colombia
colombo	colombo
colorado	colorado
colosseum	colosseum
columbia	columbia
columbus	columbus
come	come
comeback	comeback
comet	comet
cosa	cosa
costa	costa
counterstrike	counterstrike
country	country
county	county
cover	cover
craig	craig
crazy	crazy
crick	crick
cricket	cricket
criss	criss
cruz	cruz
crüe	crüe
cupen	the cup
cykel	bicycle
cykeln	cycle
cyklar	bicycles
cypern	cyprus
cyrus	cyrus
da	da
dag	day
dagar	days
dagarna	the days
dagars	day
dagbladet	daily
dagbok	diary
dagen	day
dagens	today
dagliga	daily
dagligen	daily
dagligt	daily
dags	time
dagsläget	present situation
dahlén	dahlén
dahléns	dahlén
dalar	valleys
dalarna	dalarna
dalí	dali
dam	lady
damer	ladies
dancehall	dance hall
daniel	daniel
danmark	denmark
danmarks	denmark
danny	danny
dans	dance
dansk	danish
danska	danish
danske	danish
dark	dark
darwin	darwin
darwins	darwin
das	das
data	data
dateras	dates
dator	computer
datorer	pc
datorn	computer
datorspel	computer game
datum	date
dave	dave
david	david
davis	davis
day	day
de	the
debatt	debate
debatten	debate
debatter	debates
debut	debut
debutalbum	debut
debutalbumet	debut album
debuterade	debut
december	december
decennier	decades
decennierna	decades
decenniet	decade
decennium	decade
deep	deep
define	define
definiera	define
definierade	defined
definierar	defines
definieras	defined
definierat	defined
definition	definition
definitionen	defined
definitioner	definitions
definitivt	definitely
deklarerade	declared
del	part
dela	share
delad	shared
delade	partial
delades	awarded
delar	parts
delarna	parts
delas	broken
delat	shared
delats	distributed
delen	part
delhi	delhi
delning	division
delningen	pitch
dels	partly
delstat	state
delstaten	land
delstater	states
delstaterna	states
delta	participate
deltagande	participation
deltagare	contestant
deltagarna	participants
deltagit	participated
deltar	part
deltog	participated
delvis	partly
dem	those
demens	dementia
demo	demo
demografi	demography
demografiska	demographic
demokrati	democracy
demokratier	democracies
demokratin	democratic
demokratisk	democratic
demokratiska	democratic
demokratiskt	democratic
demonstrationer	demonstrations
den	the
denna	this
denne	he
dennes	his
dennis	dennis
densamma	same
densitet	density
densiteten	density
departement	department
depolarisering	depolarization
depp	depp
depression	depression
depressionen	depression
depressioner	depression
der	where
deras	their
derivata	derivative
derivatan	derivative
derivator	derivatives
design	design
desmond	desmond
dess	its
dessa	these
dessförinnan	before
dessutom	also
desto	the
det	the
detalj	detail
detaljer	details
detroit	detroit
detsamma	the same
detta	this
deuterium	deuterium
development	development
diabetes	diabetes
diagnos	diagnosis
diagnosen	diagnosis
diagnoser	diagnoses
dialekt	dialect
dialekter	dialects
dialekterna	dialects
dialog	dialogue
diamant	diamond
diamanter	diamonds
diameter	diameter
diamond	diamond
dianno	dianno
dickens	dicken's
dickinson	dickinson
diego	diego
digerdöden	the black death
digital	digital
dikt	poem
diktator	dictator
diktatorn	dictator
diktatur	dictatorship
diktaturen	dictatorship
dikter	poetry
dillinger	dillinger
dimensioner	dimensions
din	your
dinosaurier	dinosaurs
dinosaurierna	dinosaurs
diplomatiska	diplomatic
direkt	immediately
direkta	direct
direktör	director
diskar	disks
diskografi	discography
diskriminering	discrimination
diskussion	discussion
diskussioner	discussions
diskutera	discuss
diskuterades	discussed
diskuteras	discussed
diskuterats	discussed
disney	disney
disneys	disney
distinkt	distinct
distinkta	distinct
distribution	distribution
distributioner	distributions
distrikt	district
distriktet	district
dit	there
ditt	your
dittills	thus far
diverse	some
division	division
divisionen	division
dj	dj
djup	depth
djupa	deep
djupare	deeper
djupt	deep
djur	animal
djurarter	species
djuren	animals
djurens	animals
djuret	animal
djurgården	djurgården
djurgårdens	djurgården's
djävulen	devil
dna	dna
dns	dns
dock	nevertheless
dog	died
doktor	doctor
dokument	documents
dokumenterade	documented
dokumentär	documentary
dollar	dollar
dom	judgment
domare	judge
domaren	judge
domen	judgment
dominans	dominance
dominera	dominate
dominerade	dominated
dominerades	dominated
dominerande	dominant
dominerar	dominates
domineras	dominated
dominerat	dominated
domkyrka	cathedral
domkyrkan	cathedral
domstol	court
domstolar	courts
domstolen	court
don	don
donald	donald
donau	the danube
donna	donna
dop	baptism
dopamin	dopamine
dos	dosage
dotter	daughter
dottern	daughter
downs	down
dr	dr
dra	drag
drabbade	affected
drabbades	suffered
drabbar	affecting
drabbas	affected
drabbat	affected
drabbats	affected
drag	features
dragit	preferred
drama	drama
dramat	drama
dramaten	dramatic
dramatiker	playwright
dramatiska	dramatic
dramatiskt	dramatically
dramer	dramas
draperi	curtain
drar	earn
dras	drawn
dream	dream
drev	drove
drevs	concentrated
dricka	drink
dricker	drink
drift	operation
driva	drive
drivande	driving
driver	drive
drivs	run
drog	drug
drogen	drug
droger	drugs
drogmissbruk	drug abuse, substance abuse, drug addiction
drogs	coated
drottning	queen
drottningen	queen
dryck	drink
drycken	beverage
drycker	beverages
drygt	over
dräkt	costume
dröja	take
dröjde	was not until
dröm	dream
drömmar	dreams
dsmiv	dsm-iv
du	you
dubai	dubai
dubbel	double
dubbelt	double
dubbla	double
dublin	dublin
duett	duet
dvd	dvd
dvs	i.e.
dvärg	dwarf
dvärgar	dwarves
dy	younger
dygn	day
dygnet	day
dyker	dives
dylan	dylan
dylikt	such
dynamiska	dynamic
dyrare	more expensive
dyraste	most expensive
dyrt	expensive
dä	then
däggdjur	mammal
däggdjuren	the mammals
där	where
därav	thereof
därefter	then
däremot	however
därför	therefore
däribland	among them
därifrån	from there
därigenom	thereby
därmed	thereby
därpå	thereon
därtill	thereto
därutöver	addition
därvid	thereby
då	then
dålig	bad
dåliga	bad
dåtidens	contemporary
dåvarande	then
dö	die
död	death
döda	kill
dödad	killed
dödade	killed
dödades	killed
dödar	kills
dödas	killed
dödat	killed
döden	death
dödlig	lethal
dödligheten	mortality
dödligt	deadly
dödsfall	death
dödshjälp	euthanasia
dödsoffer	death victim
dödsorsaken	cause of death
dödsstraff	death penalty
dödsstraffet	death penalty
dök	turned
dömande	judicial
dömd	convicted
dömdes	sentenced
döpt	named
döpte	baptized
döptes	named
dör	dies
dött	dead
döttrar	daughters
e	e
earl	earl
earth	earth
ebba	ebba
economic	economic
ecuador	ecuador
ed	ed
eddie	eddie
edgar	edgar
edison	edison
edith	edith
edmund	edmund
edvard	edvard
edwall	edwall
edward	edward
edwards	edward's
edwin	edwin
effekt	effect
effekten	effect
effekter	effects
effekterna	effects
effektiv	effective
effektiva	effective
effektivt	effective
efter	after
efterfrågan	demand
efterföljande	following
efterföljare	follower
efterhand	post
efterkrigstiden	the post-war period
efternamn	last name
eftersom	since
efterträdare	successor
efterträddes	succeeded
eftervärlden	posterity
efteråt	afterwards
egen	own
egendom	property
egenskap	property
egenskaper	characteristics
egenskaperna	properties
egentlig	real
egentliga	actual
egentligen	actually
eget	own
egna	own
egypten	egypt
egyptens	egypt
egyptiska	egyptian
eiffeltornet	the eiffel tower
einstein	einstein
einsteins	einstein
ej	not
eker	spoke
eklund	eklund
ekman	ekman
ekologi	ecology
ekologiska	organic
ekonomi	economy
ekonomier	economies
ekonomin	economy
ekonomisk	economic
ekonomiska	economic
ekonomiskt	economic
ekosystem	ecosystem
ekr	ad
ekvatorn	equator
eld	fire
elden	fire
electric	electric
elektricitet	electricity
elektrisk	electrical
elektriska	electric
elektriskt	electric
elektromagnetisk	electromagnetic
elektron	electron
elektroner	electrons
elektronik	electronics
element	element
eleonora	eleonora
elever	students
eleverna	the pupils
elin	elin
elisabeth	elisabeth
elit	elite
eliten	elite
elitserien	elitserien
eller	or
elton	elton
elva	eleven
elvis	elvis
em	european championship
emellan	between
emellanåt	occasionally
emellertid	however
emi	emi
emigrerade	emigrated
emil	emil
eminem	eminem
emma	emma
emmanuel	emmanuel
emo	emo
empati	empathy
empire	empire
en	one
ena	one
enade	united
enades	agreed
enastående	exceptional
enat	united
enbart	only
encyclopedia	encyclopedia
enda	only
endast	only
ende	only
energi	energy
energikälla	energy
energikällor	energy
energin	energy
energy	energy
engagemang	commitment
engagerad	engaged
engagerade	dedicated
engels	engels
engelsk	english
engelska	english
engelskan	english
engelskans	the english
engelske	english
engelskspråkiga	english
engelsmännen	english
england	england
englands	england
english	english
enhet	unit
enheten	unit
enheter	units
enhetlig	uniform
enighet	agreement
enkel	simple
enkelt	easy
enkla	easy
enklare	easier
enklaste	easiest
enlighet	according
enligt	according to
enorm	enormous
enorma	enormous
enormt	gigantic
ens	even
ensam	alone
ensamma	alone
enskild	individual
enskilda	individual
enskilt	single
enstaka	single
entertainment	entertainment
enzymer	enzymes
ep	ep
epicentrum	epicentre
epok	epoch
epoken	epoch
epost	e-mail
er	your
era	era
eran	era
erbjuda	offer
erbjuder	offers
erbjöd	offered
erbjöds	offered
erektion	erection
erfarenhet	experience
erfarenheter	experiences
erhållit	obtained
erhöll	obtained
eric	eric
ericsson	ericsson
erik	erik
eriksson	eriksson
eritrea	eritrea
erkänd	recognized
erkända	recognized
erkände	confession
erkänna	recognize
erkännande	recognition
erkänner	recognize
erkänt	recognized
ernest	ernest
ernman	ernman
ernst	ernst
eros	eros
ersatt	replaced
ersatte	replaced
ersattes	replaced
ersatts	replaced
ersätta	replace
ersättare	replacement
ersättning	replacement
ersätts	replaced
erövra	conquer
erövrade	conquered
erövrades	conquered
erövring	conquest
erövringar	conquest
erövringen	conquest
estetik	esthetics
estetiska	aesthetic
estland	estonia
estniska	estonian
et	et
etablera	establish
etablerad	established
etablerade	established
etablerades	established
etablerat	established
etanol	ethanol
etik	ethics
etiken	ethics
etiopien	ethiopia
etiopiska	ethiopian
etiska	ehtical
etnicitet	ethnicity
etnisk	ethnic
etniska	ethnic
etniskt	ethnic
ett	one
etta	one
etymologi	etymology
eu	eu
euro	euro
euron	euro
euroområdet	eurozone
europa	europe
europacupen	european cup
europaparlamentet	calls
europarådet	council of europe
europas	europe
europe	european
european	european
europeisk	european
europeiska	european
européer	europeans
européerna	europeans
eurovision	eurovision
eus	eu
eva	eva
evangelierna	the gospels
evangeliska	evangelical
evans	evans
evenemang	event
eventuell	eventual
eventuella	any
eventuellt	possibly
evert	evert
everton	everton
eviga	eternal
evigt	forever
evolution	evolution
evolutionen	evolution
evolutionsteorin	theory of evolution
ex	ex
exakt	accurately
exakta	exact
examen	exam
exempel	example
exempelvis	e.g.
exemplar	copy
exemplet	example
exil	exile
existens	existence
existensen	existence
existera	exist
existerade	existed
existerande	existing
existerar	exists
existerat	existed
exklusiv	exclusive
expandera	expand
expansion	expansion
expansionen	expansion
expedition	expedition
expeditionen	expedition
expeditioner	expeditions
experiment	experiment
experimenterade	experimented
experter	experts
explosionen	the explosion
export	export
exporten	exports
express	express
expressen	express
externa	external
extra	optional
extrem	extreme
extrema	extreme
extremt	extreme
fabriker	factories
facebook	facebook
fackföreningar	unions
facto	facto
facupen	fa cup
fader	father
fadern	father
faderns	the father's
fagocyt	phagocyte
fakta	fact
faktiska	actual
faktiskt	actually
faktor	factor
faktorer	factors
faktorn	factor
faktum	fact
fall	case
falla	fall
fallen	cases
faller	fall
fallet	case
fallit	fallen
falska	false
falskt	false
familj	family
familjen	family
familjens	family
familjer	families
familjerna	families
fan	devil
fann	found
fanns	was
fans	fans
fansen	fans
far	father
fara	danger
farbror	uncle
farfar	paternal grandfather
farlig	dangerous
farliga	dangerous
farligt	dangerous
fars	father's
fart	speed
fartyg	ship
fartyget	ship; vessel
fas	phase
fascism	fascism
fascismen	fascism
fascisterna	fascists
fascistiska	fascist
fasen	phase
faser	phases
fast	fixed
fasta	solid
fastigheter	real estates
fastlandet	mainland
fastställa	determine
fastställdes	set
fastän	although
fat	fat
fatta	take
fattas	taken
fattiga	poor
fattigare	poorer
fattigaste	poorest
fattigdom	poverty
fattigdomen	poverty
fauna	fauna
fbi	fbi
fc	fc
fci	fci
fd	ex
feber	fever
februari	february
federal	federal
federala	federal
federation	federation
federationen	federation
fel	faults
felaktig	incorrect
felaktiga	false
felaktigt	incorrect
felix	felix
fem	five
feminism	feminism
feminismen	feminism
feminister	feminists
feministiska	feminist
femte	fifth
femton	fifteen
fenomen	phenomenon
fenomenet	phenomenon
feodala	feudal
ferdinand	ferdinand
fermentering	fermentation
fernando	fernando
fest	party
fester	treats
festival	festival
festivalen	festival
festivaler	festivals
fett	fat
ff	ff
fick	got
fiende	enemy
fienden	enemy
fiender	enemies
fifa	fifa
figur	figure
figuren	figure
figurer	figures
figurerna	figures
fiktion	fiction
fiktiv	fictive
fiktiva	romantic
fil	master of
filip	filip
filippinerna	the philippines
film	film
filmatiserats	filmed
filmen	film
filmens	film
filmer	movies
filmerna	films
filmografi	filmography
filosofen	philosopher
filosofer	philosophers
filosofi	philosophy
filosofin	philosophy
filosofins	philosophy
filosofisk	philosophical
filosofiska	philosophical
fina	fine
final	final
finalen	final
finansiella	financial
finansiera	finance
finansieras	financed
finansiering	financiation
finanskrisen	financial crisis
finger	finger
fingrar	fingers
finland	finland
finlands	finland
finländska	finnish
finna	found
finnas	be
finner	finds
finns	exist
finsk	finnish
finska	finnish
fira	celebrate
firade	celebrated
firades	celebrated
firandet	celebrate
firar	celebrates
firas	celebrated
fire	fire
fisk	fish
fiskar	fish
fiske	fishing
fission	fission
fjorton	fourteen
fjädrar	spring
fjärde	fourth
fjärdedel	quarter
flagga	flag
flaggan	flag
flaggor	flags
flames	flames
flamländska	flemish
flandern	flanders
fler	more
flera	several
flertal	multiple
flertalet	most
flest	most
flesta	most
flicka	girl
flickan	girl
flickor	girls
flickvän	girlfriend
flight	rate
flitigt	actively
flod	river
floden	the river
floder	rivers
floderna	rivers
flora	flora
florens	florence
florida	florida
flotta	fleet
flottan	navy
floyd	floyd
fly	escape
flydde	escaped
flyg	flight
flyga	fly
flygande	flying
flygbolag	airline
flyger	fly
flygplan	airplane
flygplats	airport
flygplatsen	airport
flygplatser	airports
flygvapnet	air force
flykt	escape
flyktingar	refugees
flyr	flees
flytande	liquid
flyter	flows
flytt	move
flytta	move
flyttades	moved
flyttar	move
flyttas	moved
flyttat	moved
flöde	flow
flög	flew
fn	un
fns	un
fokus	focus
fokusera	focus
fokuserade	focused
fokuserar	focus
folk	people
folke	folke
folken	peoples
folket	people
folkets	people
folkgrupper	communities
folklig	popular
folkliga	folk
folkmord	genocide
folkmordet	genocide
folkmun	popularly
folkmusik	folk music
folkmängd	population
folkmängden	population
folkomröstning	referendum
folkpartiet	peoples party
folkrepubliken	people's republic
folkrikaste	populous
folkräkning	census
folkräkningen	census
folkslag	peoples
folktro	folklore
folkvalda	elected
fontsizes	fontsizes
football	football
force	force
ford	ford
fordon	vehicle
form	form
format	format
formatet	format
formel	formula
formell	formal
formella	formal
formellt	formally
formen	form
former	forms
formerna	forms
forna	former
fornnordiska	norse
forntida	ancient
forsberg	forsberg
forskare	researcher
forskaren	researcher
forskarna	scientists
forskning	research
forskningen	research
fort	fast
fortfarande	still
fortplantning	reproduction
fortsatt	continued
fortsatta	further
fortsatte	continued
fortsätta	continue
fortsätter	continues
fortsättning	continuation
fortsättningen	continue
forum	forum
fossil	fossil
fossila	fossil
foster	fetal
fot	foot
fotbeklädnad	footwear
fotboll	football
fotbollen	football
fotbollslandslag	football team
fotbollsspelare	footballers
foten	foot
fotnoter	footnotes
foto	photo
fotografier	photographs
foton	photos
fotosyntesen	photosynthesis
fragment	fragment
fralagen	the fra law
fram	front
framför	in front of
framföra	present
framförallt	especially
framförde	performed
framfördes	expressed
framförs	expressed
framfört	forward
framförts	forward
framgång	success
framgångar	successes
framgångarna	successes
framgången	success
framgångsrik	successful
framgångsrika	successful
framgångsrikt	successfully
framgår	clear
framsteg	progress
framställa	produce
framställning	production
framställs	prepared
framstående	prominent
framtid	future
framtida	future
framtiden	the future
framträdande	prominent
framträdanden	performance
framträdde	appeared
framträder	stand
framåt	forward
francis	francis
francisco	fransisco
franco	franco
franklin	franklin
frankrike	france
frankrikes	france
fransk	french
franska	french
franske	french
franskt	french
fransmännen	french
franz	franz
français	francais
fred	peace
freddie	freddie
freddy	freddy
freden	peace
fredliga	peaceful
fredrik	fredrik
fredsbevarande	peace
fredspris	prize
fredspriset	peace prize
freedom	freedom
freja	joe
frekvens	frequency
freud	freud
fri	free
fria	free
friedrich	friedrich
frigörelse	liberation
frigörs	released
frihet	freedom
friheten	freedom
frihetliga	libertarian
friidrott	athletics
frisk	healthy
friska	healthy
fristående	independent
fritid	free time
fritt	free
fritz	fritz
frivillig	voluntary
frivilliga	voluntary
frivilligt	voluntary
frodo	frodo
from	from
front	front
fronten	front
fru	wife
frukt	fruit
fruktade	feared
frälsning	salvation
främja	promote
främmande	foreign
främre	front
främst	foremost; primarily; chiefly
främsta	primary
främste	chief
fråga	question
frågade	asked
frågan	the question
frågor	issues
frågorna	issues
från	from
frånträde	withdrawal
frånvaro	absence
fröken	miss
fröväxter	seed plants
fss	fss
fuglesang	fuglesang
fuktiga	damply
fuktigt	moist
full	full
fulla	full
fullständig	full
fullständiga	full
fullständigt	completely
fullt	full; fully; completely
fungera	work
fungerade	did
fungerande	functioning
fungerar	functions
funktion	feature
funktionella	functional
funktionen	function
funktioner	functions
funktionerna	functions
funnit	found
funnits	found
fursten	prince
fusion	fusion
fusionen	the fusion
futharkens	futhark
fylla	fill
fyllde	filled
fyller	turns
fynd	finding; finds
fynden	finds
fyra	four
fyrtio	forty
fysik	physics
fysikaliska	physical
fysiker	physicist
fysiologi	physiology
fysiologiska	physiological
fysisk	physical
fysiska	physical
fysiskt	physically
fält	field
fältet	the field
fälttåg	campaign
fängelse	prison
fängelsestraff	imprisonment
fängelset	prison
fängslade	imprisoned
fängslades	imprisoned
färdas	travel
färdig	finished
färdiga	actual
färg	color
färgade	colored
färgen	color
färger	colors
färgerna	colors
färre	less
färöarna	faroe islands
fäste	attachment
fästning	fortress
få	get
fåfotingar	pauropoda
fågel	bird
fågelarter	species
fågelhundar	bird dogs
fåglar	birds
fåglarna	the birds
fåglarnas	birds
fånga	capture
fångar	prisoners
fångenskap	captivity
får	may
fåtal	few
fått	got
föda	food
född	born
födda	born
födde	gave birth too
föddes	born
födelse	birth
födelsedag	birthday
födelsetal	birth
föder	give birth of
föds	born
födseln	birth
föga	little
följa	follow
följaktligen	consequently
följande	following
följas	followed
följd	sequence
följde	followed
följden	sequence
följder	impact
följdes	followed
följer	resulting
följeslagare	companion
följs	followed
följt	followed
föll	fell
fönster	window
för	for
föra	bring
föranledde	brought about
föras	be
förband	units; formations; bound (themselves)
förbi	past
förbindelse	connection
förbindelser	relations
förbinder	connects
förbjuda	ban
förbjuden	prohibited
förbjuder	prohibiting
förbjudet	prohibited
förbjudna	forbidden
förbjöd	forbid
förbjöds	forbidden
förblev	remained
förblir	remains
förbränning	combustion
förbud	prohibition
förbudet	prohibition
förbund	union
förbundet	association
förbundskapten	coach
förbundsrepubliken	federal republic
förbundsstat	federal state
förbättra	improve
förbättrade	improved
förbättringar	improvement
förde	brought
fördel	advantage
fördelade	distributed
fördelar	advantages
fördelas	distributed
fördelen	advantage
fördelning	distribution
fördelningen	distribution
fördes	sea were entered
fördomar	bias
fördrag	treaty
fördragen	treaties
fördraget	treaty
fördrevs	was banished
före	before
förebild	role model
förebyggande	preventing
föredrar	prefer
föredrog	preferred
förefaller	appears
föregående	previous
föregångare	predecessor
föregångaren	predecessor
förekom	occurred
förekomma	occur
förekommande	occuring
förekommer	present
förekommit	occurred
förekomst	presence
förekomsten	presence
föreligger	exists
föremål	subject
förena	combine
förenade	joined
förening	association
föreningar	associations
föreningen	association
förenklat	simplified
förenta	united
föreslagit	proposed
föreslagits	suggested
föreslog	suggested
föreslogs	proposed
föreslår	suggest
förespråkade	advocated
förespråkar	advocate
förespråkare	advocate
föreställa	imagine
föreställande	depicting
föreställer	represents
föreställning	show
föreställningar	performances
föreställningen	show
företag	business
företagen	companies
företaget	now
företagets	company
företeelse	phenomenon
företeelser	phenomena
företrädare	representatives
företräder	represents
författare	author
författaren	author
författarna	writers
författarskap	authorship
författning	constitution
författningen	constitution
förfäder	ancestors
förföljelse	persecution
förföljelser	persecution
förgäves	in vain
förhandla	negotiate
förhandlingar	negotiations
förhandlingarna	negotiations
förhindra	prevent
förhindrar	prevent
förhistoria	prehistory
förhistorisk	prehistoric
förhärskande	predominant
förhållande	relationship
förhållanden	conditions
förhållandena	conditions
förhållandet	ratio
förhållandevis	relatively
förhåller	relationship
förhöjd	enhanced
förintelsen	the genocide
förklara	explain
förklarade	explained
förklarades	declared
förklaras	explained
förklarat	explained
förklaring	explanation
förklaringar	explanations
förklaringen	the explanation
förknippad	associated
förknippade	associated
förknippas	associated
förkortas	shortened
förkortat	abbreviated
förkortning	abbreviation
förkortningar	abbreviations
förlag	magazine
förlaget	publisher
förlopp	course
förlora	lose
förlorade	lost
förlorades	lost
förlorar	loses
förlorat	lost
förlust	loss
förlusten	loss
förluster	loss
förlusterna	losses
förlängning	extension
förlängningen	extension
förmedla	pass; express; mediate
förmodligen	probably
förmåga	ability
förmågan	the ability
förmågor	abilities
förmån	benefit
förmögenhet	fortune
förnuft	sense
förnuftet	sense
förorter	suburbs
förr	before
förra	last
förrän	before
förs	out
församling	assembly
församlingar	assemblies
församlingen	assembly
förslag	proposal
förslaget	proposal
först	first
första	first
förstaplatsen	first place
förste	first
förstnämnda	first
förstod	understood
förstärka	strengthen
förstå	understand
förståelse	understanding
förståelsen	understanding
förstår	understand
förstås	course
förstöra	destroy
förstördes	was destroyed
förstörelse	destruction
försvann	disappeared
försvar	defense
försvara	defend
försvarade	defended
försvarare	defender
försvaret	defense
försvarets	defense
försvarsmakt	armed
försvarsmakten	defense
försvarsminister	defense
försvinna	disappear
försvinner	disappear
försvunnit	disappeared
försäkra	make sure
försäljning	sale
försäljningen	sales
försämrades	worsened
försök	attempt
försöka	try
försöken	attempts
försöker	trying
försökt	tried
försökte	tried
försörja	support
försörjde	supported
försörjning	sustention
fört	pre
förteckning	list
förtjust	fond
förtroende	trust
förtryck	opression
förts	transferred
förut	before
förutom	except
förutsätter	requires
förutsättning	provided
förutsättningar	conditions
förutsättningarna	conditions
förvaltning	management
förvaras	stored
förväntade	expected
förväntas	expected
förväntningar	expectations
förväxla	mistake
förväxlas	confused
föräldrar	parents
föräldrarna	the parents
förälskad	in love
förändra	change
förändrade	changed
förändrades	changed
förändras	change
förändrats	changed
förändring	change
förändringar	changes
förändringarna	changes
förändringen	change
förödande	devastating
fötter	feet
fötterna	feet
fötts	born
führer	fuhrer
gabriel	gabriel
gaga	gaga
galax	galaxy
galaxer	galaxies
galilei	galilei
galileo	galileo
gallagher	gallagher
galleri	gallery
gallien	gaul
gamla	old
gamle	old
gammal	old
gammalt	old
gandalf	gandalf
gandhi	gandhi
gandhis	gandhi
ganska	quite
garantera	guarantee
garanterar	ensures
garvey	garvey
gary	gary
gas	gas
gasen	gas
gata	street
gatan	street
gates	gates
gator	streets
gatorna	streets
gav	gave
gavs	was given
gaza	gaza
gazaremsan	gaza strip
ge	give
gemensam	common
gemensamma	common
gemensamt	commonly
gemenskap	community
gemenskapen	community
gemenskaperna	communities
gen	gene
genast	immediately
genen	gene
gener	genes
general	general
generalen	general
generalguvernören	governor general
generalsekreterare	secretary general
generation	generation
generationen	generation
generationer	generations
generell	general
generella	general
generellt	generally
generna	genes
genetik	genetics
genetisk	genetic
genetiska	genetic
genetiskt	genetically
genom	by
genombrott	breakthrough
genombrottet	breakthrough
genomför	carry
genomföra	implement
genomföras	performed
genomförde	performed
genomfördes	was
genomförs	performed
genomfört	completed
genomförts	out
genomgick	underwent
genomgripande	good
genomgående	through
genomgår	undergoing
genomgått	passed
genomslag	impact
genomsnitt	average
genomsnittet	average
genomsnittlig	average
genomsnittliga	average
genre	genre
genren	genre
genrer	genres
gentemot	against
genus	gender
geografi	geography
geografisk	geographical
geografiska	geographic
geografiskt	geographically
geologi	geology
geologiska	geological
geologiskt	geological
geomorfologi	geomorphology
georg	georgian
george	george
georges	georges
georgien	georgia
georgier	georgian
ger	gives
germanska	germanic
ges	given
gestalt	figure
gestalter	figures
gett	given
ghana	ghana
gia	gia
gick	went
gift	married
gifta	married
gifte	married
gifter	marries
giftermål	marriage
giftsnokar	elapidae
gigantiska	gigantic
gillade	liked
gillar	like
giovanni	giovanni
girl	girl
girls	girls
gisslan	hostage
gitarr	guitar
gitarrist	guitarist
gitarristen	guitarist
givaren	donor
given	given
givet	given
givetvis	naturally
givit	given
givits	given
gjord	made
gjorda	made
gjorde	did
gjordes	was
gjort	done
gjorts	done
glad	happy
glada	happy
glas	glass
glenn	glenn
global	global
globala	global
globalt	global
globe	globe
globen	the globe
gloria	gloria
glukos	glucose
glädje	joy
glödlampor	lightbulbs
go	go
god	good
goda	good
godkände	approved
godkändes	approved
godkänna	approve
godkännande	approval
godkännas	approved
godkänt	approved
gods	goods
goebbels	geobbels
gogh	gogh
golf	golf
golvet	the floor
gom	palate
google	google
gorbatjov	gorbachev
gordon	gordon
got	got
gotiska	gothic
gotland	gotland
gotlands	gotland
gott	good
grace	grace
grad	grade
graden	rate
grader	degrees
gradvis	gradually
grafit	graphite
graham	graham
grammatik	grammar
grammis	grammy
grammy	grammy
gran	spruce
grand	grand
grande	grand
grannar	neighbors
granne	neighbour
grannlandet	the neighbouring country
grannländer	neighboring countries
grannländerna	neighbors
granska	review
granskning	review
grant	grant
gratis	free
grav	grave
graven	grave
gravid	pregnant
graviditet	pregnancy
graviditeten	pregnancy
gravitation	gravitation
gray	gray
greker	greeks
grekerna	greeks
grekisk	greek
grekiska	greek
grekiskans	greek
grekland	greece
greklands	greece
gren	branch
grenar	branches
grenen	branch
greps	was arrested
greve	count
griffin	griffin
griffon	griffon
grovt	rough
grund	"in the context: ""på grund"" = because of"
grunda	base
grundad	based
grundade	founded
grundades	founded
grundande	founding
grundandet	founding
grundar	found
grundare	founder
grundaren	founder
grundarna	founders
grundas	based
grundat	founded
grunden	basis
grunder	bases
grundlag	constitution
grundlagen	constitution
grundläggande	primary
grundskolan	elementary school
grundämne	element
grundämnen	elements
grundämnet	element
grupp	group
gruppen	group
gruppens	group
grupper	groups
grupperingar	groupings
grupperna	groups
gruppspelet	groupplay
gräns	limit
gränsar	border
gränsen	limit
gränser	limits
gränserna	border
gräs	grass
gräslök	chive
grå	gray
grön	green
gröna	green
grönland	greenland
grönsaker	vegetables
grönt	green
grönwall	grönwall
guatemala	guatemala
gud	god
gudar	gods
gudarna	gods
gudarnas	gods
guden	god
gudinnan	the godess
gudom	deity
gudomlig	divine
gudomliga	divine
guds	god
guevara	guevara
guide	guide
guillou	guillou
guinea	guinea
gul	yellow
gula	yellow
guld	gold
guldbollen	golden ball
gunnar	gunnar
guns	guns
gunwer	gunwer
gustaf	gustaf
gustafs	gustaf
gustafsson	gustafsson
gustav	gustav
gustavs	gustav
guvernör	governor
guyana	guyana
gyllene	golden
gymnasiet	high school
gymnasium	gymnasium
gälla	be valid
gällande	current
gällde	applied
gäller	of
gäng	group
gänget	the group
gärna	i'd love to
gärning	act
gärningar	works
gärningsmannen	perpetrator; offender
gäst	guest
gäster	guests
gävle	gävle
gå	go
gång	time
gången	time
gånger	times
gångna	past
går	goes
gård	farm
gården	farm
gått	gone
gåva	gift
gör	makes
göra	do
göran	göran
göras	done
göring	attachment
görs	is
gösta	gösta
göta	göta
götaland	götaland
göteborg	gothenburg
göteborgs	gothenburg
h	h
ha	have
haag	the hague
haber	haber
haddock	haddock
hade	had
haft	had
haile	haile
haiti	haiti
hall	hall
halland	halland
halloween	halloween
hallucinationer	hallucinations
halmstad	halmstad's
halmstads	halmstad's
hals	throat
halsen	throat
halt	stop; level
halv	half
halva	half
halvan	half
halvklotet	hemisphere
halvt	half
halvön	the peninsula
hamas	hamas
hamburg	hamburger
hamilton	hamilton
hamlet	hamlet
hammarby	hammarby
hamn	port
hamna	end
hamnade	ended
hamnar	ports
hamnat	got
hamnen	port
hampa	hemp
han	he
hanar	males
hand	hand
handboll	handball
handel	trade
handeln	trade
handels	trade
handelsmän	merchants
handelspartner	trading partner
handen	hand
handla	act
handlade	was
handlande	act
handlar	deal
handling	action
handlingar	actions
handlingen	act
hanen	male
hanhon	he/she
hann	could
hannah	hannah
hannar	males
hans	his
hansson	hansson
hantera	manage
hantverk	crafting
hantverkare	craftsman
har	has
harald	harald
harris	harris
harrison	harrison
harry	harry
hasch	hashish
hastighet	speed
hastigt	rapidly
hat	hatred
hatar	hate
hav	sea
have	have
haven	the seas
havet	sea
havets	sea
havs	at sea
havskattfiskar	catfishes
havsnivån	sea level
hawaii	hawaii
hawking	hawking
hc	h.c.
hdmi	hdmi
he	he
heart	heart
heath	heath
heaven	heaven
hebreiska	hebrew
hedersdoktor	honorary doctor
hegel	hegel
heinrich	heinrich
heinz	heinz
hel	whole
hela	whole
helena	helena
helgdagar	holidays
helhet	whole
helig	holy
heliga	holy
helige	holy
heligt	holy
helium	helium
hell	hell
heller	either
hellre	rather
hells	hell
hellström	hellström
helsingborg	helsingborg
helsingborgs	helsingborg
helsingfors	helsinki
helsingör	helsingor
helst	anyone
helt	completely
helvetet	hell
hem	home
hemingway	hemingway
hemland	homeland
hemlandet	homeland
hemlig	secret
hemliga	secret
hemlighet	secret
hemligt	secret
hemma	home
hemmaarena	home ground
hemmaplan	home
hemmet	home
hemsida	website
hendrix	hendrix
henne	her
hennes	her
henri	henri
henrik	henrik
henriks	henry
henry	henry
hepatit	hepatite
herbert	herbert
hercegovina	herzegovina
hergé	hergé
heritage	heritage
herman	herman
hermann	hermann
heroin	heroin
herr	mister
herrar	men
herre	lord
herren	lord
herrens	lord
herrlandskamper	men's international contest
herrlandslag	football team
hertig	duke
het	hot
heta	hot
heter	called
hett	hot
hette	named
hexadecimalt	hexa-decimal
heydrich	heydrich
high	high
himlakroppar	celestial bodies
himlen	heaven
himmel	sky
himmler	himmler
himmlers	himmler
hinder	obstacle
hindra	prevent
hindrade	prevented
hindrar	prevent
hindu	hindu
hinduer	hindu
hinduiska	hindu
hinduism	hinduism
hinduismen	hindu
hinner	have time to
hiroshima	hiroshima
his	his
hisingen	hisingen
historia	history
historien	history
historiens	history
historier	stories
historik	history
historiker	historian
historikern	historian
historisk	historical
historiska	historical
historiskt	historic
history	history
hit	here
hitler	hitler
hitlers	hitler
hits	hits
hitta	see
hittade	found
hittades	found
hittar	finds
hittas	be found
hittat	found
hittats	found
hittills	date
hiv	hiv
hjalmar	hjalmar
hjälp	help
hjälpa	help
hjälper	help
hjälpmedel	aid
hjälpt	helped
hjälpte	helped
hjärna	brain
hjärnan	brain
hjärnans	brain
hjärta	heart
hjärtat	heart
hms	hms
ho	ho
hockey	hockey
holland	holland
hollywood	hollywood
holländska	dutch
holm	holm
homo	homo
homogen	homogenous
homosexualitet	homosexuality
homosexuell	homosexual
homosexuella	homosexual
hon	she
honan	female
honom	him
honor	ära
hopp	hope
hoppa	skip
hoppade	jumped
hoppades	hoped
hoppas	hope
hormoner	hormons
horn	horn
hos	at
hotad	threatened
hotade	threatened
hotar	threatens
hotel	hotel
hotell	hotel
hotellet	hotel
hotet	the threat
house	house
houston	houston
hov	court
hovet	court
hovrätten	the court of appeal
how	how
howard	howard
hud	skin
huden	skin
hudfärg	color
hughes	hughes
hugo	hugo
human	human
humanism	humanism
humanismen	humanism
humanistiska	humane
humle	hop
humor	humour
humör	temper
hund	dog
hundar	dogs
hunden	the dog
hundra	hundred
hundraser	alternative strains
hundratal	hundred
hundratals	hundreds
hundratusentals	hundreds of thousands
hunnit	reached
hur	how
huruvida	whether
hus	house
husen	houses
huset	house
hushåll	household
huskvarna	huskvarna
hussein	hussein
hustru	wife
hustrun	wife
huvud	head
huvudartikel	main article
huvuddelen	main part
huvudet	head
huvudkontor	central office
huvudort	capital
huvudperson	main character
huvudrollen	the main role
huvudsak	substantially
huvudsakliga	main
huvudsakligen	generally
huvudstad	capital
huvudstaden	capital
huvudstäder	capitals
huvudvärk	headache
huxley	huxley
hyllade	celebrated
hyllning	tribute; homage
hypotes	hypothesis
hypotesen	hypothesis
hypoteser	hypotheses
hyser	has
häcklöpning	hurdles
hälft	half
hälften	half
hällristning	petroglyph
hälsa	tell (him i said hi)
hämnd	revenge
hämta	retrieve
hämtade	brought
hämtar	download
hämtat	collected
hända	happen
hände	happened
händelse	event
händelsehorisonten	event horizon
händelsen	event
händelser	handelsar
händelserna	the events
händer	happens
händerna	hands
hänga	hang
hänger	bag
hänsyn	regard
hänt	happened
hänvisa	refer
hänvisade	referred
hänvisar	refers
hänvisning	reference
här	here
härifrån	from here
härkomst	origin
härledas	derived
härrör	derived
härskare	ruler
härstamma	originate
härstammar	derived
härstamning	origin
häst	horse
hästar	horses
hästen	horse
hästens	horse
hävda	claim
hävdade	claimed
hävdar	assert
hävdat	claimed
håkan	chin
håkansson	hakansson
hål	hole
hålet	hole
håll	hold
hålla	keep
hållas	be
håller	holds
hållet	direction
hållit	stayed
hållning	position
hålls	held
hår	hair
hård	hard
hårda	hard
hårdare	harder
hårdast	the most
hårdrock	metal
hårdrocken	hard rock
hårdvara	hardware
håret	hair
hårt	hard
höftledsgrop	acetabulum
hög	high
höga	high
höger	right
högkvarter	headquarters
höglandet	highlands
högra	right
högre	higher
högskola	college
högskolan	science
högskolor	colleges
högst	highest
högsta	highest
högste	chief
högt	high
högtid	festival
högtider	holidays
högtryck	high pressure
höja	raise
höjd	height
höjder	heights
höjdes	increased
höjdpunkt	peak
höjer	increases
höll	hold
hölls	was
hör	hear
höra	hear
hörde	heard
hörn	corner
hörs	heard
hört	heard
höst	fall
hösten	autumn
i	in
ian	ian
iberiska	iberian
ibland	sometimes
ibm	ibm
ibn	ibn
ibrahimović	ibrahimovic
icd	icd
icke	non
ida	ida
idag	today
ideal	ideal
identifiera	identification
identifierade	identified
identisk	identical
identitet	identity
ideologi	ideology
ideologier	ideologies
ideologin	ideology
ideologiska	ideology
ideologiskt	ideology
idol	idol
idrott	sports
idéer	ideas
idén	idea
ifall	if
ifk	ifk
ifråga	in question
ifrågasatt	questioned
ifrågasatts	is questioned
ifrån	from
igelkott	hedgehog
igelkottar	hedgehogs
igelkotten	hedgehog
igelkottens	hedgehog
igen	again
igenom	through
igång	started
ihop	together
ihåg	remember
iii	iii
iiis	iii's
iis	ii's
ikea	ikea
ikon	icon
illa	bad
illegal	illegal
illegala	illegal
illinois	illinois
illuminati	illuminati
ilska	anger
image	image
imf	imf
immigranter	immigrants
immunförsvar	immune
imperiet	empire
imperium	empire
import	import
in	in
inblandad	involved
inblandade	involved
inblandning	involvement
inbördes	intermutual
inbördeskrig	civil war
inbördeskriget	civil war
indelad	divided
indelade	divided
indelas	split
indelat	divided
indelning	division
indelningar	divisions
indelningen	division
independence	independence
index	index
indian	indian
indiana	indiana
indianer	native
indianerna	indians
indianska	indian
indien	india
indiens	india
indier	indian
indierna	indians
indikerar	indicates
indirekt	indirectly
indisk	indian
indiska	indian
individ	individual
individen	individual
individens	individual
individer	individuals
individerna	individuals
individuella	individual
indoeuropeiska	indo-european
indonesien	indonesia
indonesiska	indonesian
industri	industry
industrialiserade	industrialized
industrialisering	industrialization
industrialiseringen	industrialization
industriell	industrial
industriella	industrial
industriellt	industrial
industrier	industries
industrin	industry
infaller	incident
infektion	infection
infektioner	infections
inflation	inflation
inflationen	inflation
influensa	influenza
influensan	flu
influensavirus	flu virus
influenser	influence
influerad	influenced
influerat	influenced
inflytande	influence
inflytandet	influence
inflytelserika	influential
information	information
informationen	information
infrastruktur	infrastructure
infrastrukturen	infrastructure
infödda	natives
inför	before
införa	introduce
införande	introduction
införandet	introduction
införde	introduced
infördes	introduced
infört	introduced
införts	introduced
inga	no
ingen	no
ingenjör	engineer
ingenting	nothing
inget	nothing
ingick	part
ingmar	ingmar
ingredienser	ingredients
ingrid	ingrid
ingripa	interfere
ingripande	intervention
ingvar	ingvar
ingå	part
ingående	enter into
ingår	included
ingått	concluded
inhemsk	domestic
inhemska	native
initiativ	initiative
inkluderade	included
inkluderar	include
inkluderas	included
inkluderat	including
inklusive	including
inkomst	income
inkomster	income
inkomsterna	revenue
inkomstkälla	was added to cold
inlandet	inland
inleda	initiate
inledande	initial
inledde	initiated
inleddes	initiated
inleder	initiates
inledning	introduction
inledningen	introduction
inledningsvis	initially
inleds	initiated
inlett	initiated
inletts	initiated
inlägg	post
inlärning	learning
innan	before
innanför	inside
inne	in
innebandy	floorball
innebar	meant
inneburit	meant
innebär	means
innebära	means
innebörd	meaning
innebörden	meaning
innefattar	includes
innehade	held
innehar	hold
innehas	held
innehav	owning
innehåll	content
innehålla	contain
innehållande	including
innehåller	contains
innehållet	content
innehöll	include
innersta	inner
innerstaden	inner city
inom	within
inre	internal
inrikes	domestic
inriktad	oriented
inriktade	oriented
inriktning	alignment
inriktningar	direction
inrättades	up
insats	insert
insatser	action
insekter	insects
inser	realizes
insikt	insight
inslag	element
inspelad	recorded
inspelning	recording
inspelningar	recordings
inspelningarna	recordings
inspelningen	recording
inspiration	inspiration
inspirerad	inspired
inspirerade	inspired
inspirerades	inspired
inspirerat	inspired
instabil	unstable
installera	install
instiftade	created
institut	institution
institutet	institute
institutioner	institutions
institutionerna	institutions
instruktioner	instructions
instrument	intrument
inställning	attitude
insulin	insulin
insåg	realized
inta	taken
intag	intake
inte	not
integration	integration
integritet	integrity
intellektuella	intellectual
intensiv	intensive
intensiva	intensive
intensivt	intensive
inter	inter
interaktion	interaction
interna	internal
international	international
internationell	international
internationella	international
internationellt	internationally
internet	internet
interstellära	interstellar
intervju	interview
intervjuer	interviews
intet	no
intill	next to
intog	took
intogs	was taken
intressant	interesting
intressanta	interesting
intresse	interest
intressen	interests
intresserad	interested
intresserade	interested
intresset	interest
introducerade	introduced
introducerades	introduced
intryck	impression
inträde	entry
inträffade	occurred
inträffar	occur
intäkter	income
intäkterna	the revenues
intåg	entry
inuti	inside
invadera	invade
invaderade	invaded
invaldes	elected
invandrade	immigrant
invandrare	immigrant
invandring	immigration
invasion	invasion
invasionen	invasion
inverkan	impact
investeringar	investments
invigdes	was opened
invigningen	opening
invånare	inhabitants
invånarna	residents
inåt	inwards
ip	ip
irak	iraq
irakiska	iraqi
irakkriget	iraq war
iraks	iraq
iran	iran
irans	iran's
iranska	iranian
irland	ireland
irländska	irish
isberg	iceberg
isbn	isbn
isen	ice
ishockey	ice hockey
ishockeyspelare	hockey players
islam	islam
islamisk	islamic
islamiska	islamic
islamistiska	islamic
islams	islam
island	icelandic
isländska	icelandic
iso	iso
isolerad	isolated
isolerade	isolated
isolering	isolation
isotoper	isotopes
israel	israel
israelisk	israeli
israeliska	israeli
israels	israel
istanbul	istanbul
istiden	ice age
istället	instead
isär	apart
italien	italy
italiens	italy
italiensk	italian
italienska	italian
iu	iu
ivan	ivan
ivar	ivar
iväg	away
ix	4
ja	yes
jack	jack
jackie	jackie
jackson	jackson
jacksons	jackson
jacob	jacob
jacques	jacques
jag	i
jaga	hunt
jagar	hunting
jah	jah
jakob	jacob
jakt	hunting
jakten	hunt
jamaica	jamaica
jamaicanska	jamaican
jamaicas	jamaica
james	james
jan	jan
janeiro	janeiro
januari	january
janukovytj	janukovytj
japan	japanese
japanerna	japanese
japans	japan
japansk	japanese
japanska	japanese
jarl	jarl
jason	jason
java	java
jazz	jazz
jean	jean
jeff	jeff
jefferson	jefferson
jehovas	jehovas
jennifer	jennifer
jenny	jenny
jens	jens
jensen	jensen
jersey	jersey
jerusalem	jerusalem
jerusalems	jerusalem
jesu	jesus
jesus	jesus
jihad	jihad
jim	jim
jimi	jimi
jimmy	jimmy
joachim	joachim
joakim	joakim
joan	joan
jobb	job
jobba	work
jobbade	worked
jobbar	work
jobbet	work
joe	joe
joel	joel
joey	joey
johann	johann
johannes	johannes
johans	johan's
johansson	johansson
johanssons	johansson
john	john
johnny	johnny
johnson	johnson
joker	joker
jolie	jolie
jon	jon
jonas	jonas
jonatan	jonathan
jonathan	jonathan
jones	jones
jonsson	jonsson
jord	soil
jordanien	jordan
jordbruk	agriculture
jordbruket	agricultural
jordbävning	earthquake
jordbävningar	earthquakes
jordbävningen	earthquake
jorden	earth
jordens	earth
jorderosion	earth erosion
jordskorpan	earth crust
jordytan	earth's surface
jorge	jorge
josef	joseph
joseph	joseph
josé	jose
journal	journal
journalist	journalist
journalisten	journalist
journalister	journalists
jr	junior
ju	the
juan	juan
judar	jews
judarna	jews
judarnas	jews
judas	judas
jude	jew
judendom	judaism
judendomen	the judaism
judisk	jew
judiska	jewish
judy	judy
jugoslavien	yugoslavia
jugoslaviska	jugoslavian
jul	christmas
julafton	christmas eve
juldagen	christmas day
julen	christmas
jules	jules
juli	july
julia	julia
julian	julian
julie	julie
julius	julius
juni	june
junior	junior
jupiter	jupiter
jupiters	jupiter
juridik	law
juridisk	legal
juridiska	legal
juridiskt	legally
juryn	the jury
juryns	the jury's
jussi	jussi
just	just
justice	justice
juventus	juventus
jämför	compare
jämföra	compare
jämföras	comparable
jämförelse	comparison
jämförelser	comparison
jämförelsevis	comparatively
jämfört	compared
jämlikhet	equality
jämna	even
jämnt	level
jämte	next (to)
järn	iron
järnmalm	iron ore
järnväg	railway
järnvägar	railways
järnvägarna	railways
järnvägen	railway
järnvägsnätet	rail
jönköping	jönköping
jönköpings	new
jönsson	jönsson
jönssonligan	jönssonligan
kaffe	coffee
kaffet	coffee
kairo	cairo
kalender	calendar
kalendern	calendar
kalifornien	california
kalksten	limestone
kall	cold
kalla	call
kallad	called
kallade	called
kallades	called
kallar	call
kallare	colder
kallas	called
kallat	called
kallats	called
kallblod	cold blood
kalle	kalle
kallt	cold
kalmar	kalmar
kammare	chamber
kammaren	chamber
kamp	struggle
kampanil	campanile
kampanj	campaign
kampanjen	campaign
kampen	fight
kampf	kampf
kamprad	kamprad
kan	can
kanada	canada
kanadas	canadian
kanadensiska	canadian
kanal	channel
kanalen	channel
kanaler	channels
kanarieöarna	canary islands
kandidat	candidate
kandidater	candidates
kanske	may
kant	edge
kantoner	cantons
kantonerna	cantons
kaos	chaos
kap	cape
kapacitet	capacity
kapital	capital
kapitalet	capital
kapitalism	capitalism
kapitalismen	capitalism
kapitalismens	capitalism
kapitalistiska	capitalist
kapitel	chapter
kapitulation	capitulation
kapitulerade	surrendered
kapten	captain
karakteristiska	characteristic
karaktär	character
karaktären	character
karaktärer	characters
karaktäriseras	characterized
kardinal	cardinal
karibiska	caribbean
karin	karin
karl	charles
karlsson	karlsson
karlstad	phoenix
karlstads	karlstad
karma	karma
karolinska	karolinska (institute for medicine)
karriär	career
karriären	career
karta	map
kartan	map
kartor	maps
kaspiska	caspian
kasta	throw
kastar	throws
katalanska	catalan
katalonien	catalonia
katastrofen	catastrophy
katastrofer	disasters
kate	kate
kategori	category
kategoriasiens	category of asia
kategoribrittiska	category: british
kategorier	categories
kategorieuropas	category europe
kategorifiktiva	category fictitious
kategorifödda	category: born
kategorikrigsåret	category war years
kategorikvinnor	category women
kategoriledamöter	category: members
kategorimusik	category music
kategorimän	category: men
kategorin	category
kategoriorter	category visited
kategoripersoner	category of persons
kategorirock	category:rock
kategorispelare	category player
kategorisvenska	category: swedish
kategorisvenskar	category swedes
kategorityska	category: german
katekes	catechism
katla	"katla (fictive dragon in the classic ""bröderna lejonhjärta"")"
katolicismen	catholic
katoliker	catholic
katolsk	catholic
katolska	catholic
katt	cat
kattdjur	cat
katten	the cat
katter	cats
kazakstan	kazakhstan
kedja	chain
kedjan	chain
kedjor	chains
keith	keith
kejsar	imperial
kejsardömet	empire
kejsare	emperor
kejsaren	emperor
kejsarens	emperor
kejserliga	imperial
keltiska	celtic
kemi	chemistry
kemikalier	chemicals
kemisk	chemical
kemiska	chemical
kemiskt	chemically
ken	ken
kennedy	kennedy
kenneth	kenneth
kenny	kenny
kent	kent
kenya	kenya
keramik	ceramics
kevin	kevin
kids	kids
kiev	kiev
kill	kill
kille	guy
kilometer	kilometer
kim	kim
kina	china
kinas	chinas
kinesisk	chinese
kinesiska	chinese
kings	kings
kingston	kingston
kirsten	kirsten
kiss	kiss
kjell	kjell
kl	at
klan	clan
klar	clear
klara	done
klarade	passed
klarar	pass
klart	clear
klass	grade; class
klassas	classified
klassen	the class
klasser	classes
klassificera	classifying
klassificeras	classified
klassificering	classification
klassiker	classic
klassisk	classic
klassiska	classic
klassiskt	classic
klaviatur	keyboard
klimat	climate
klimatet	environment
klimatologi	climatology
klippa	cut
klippiga	rocky
klitoris	clitoris
klockan	bell
klorofyll	cholophyll
kloster	monastery
klp	klp
klubb	club
klubbar	clubs
klubbarna	clubs
klubben	club
klubbens	club
klubblag	club
klädd	clothed
kläder	clothes
klädsel	cover
km	kilometers
km²	km²
knapp	scarce
knappast	hardly
knappt	hardly
knight	knight
knut	knot
knuten	tied to
knutna	associated
knutpunkt	hub
knutsson	knutsson
knyta	tie
knä	knee
knäppupp	knäppup
ko	cow
koalition	coalition
koden	the code
koenigsegg	koenigsegg
koffein	caffein
kognitiv	cognitive
kognitiva	cognitive
kokain	cocaine
kokpunkt	boiling point
kol	coal; charcoal
koldioxid	co
kolhydrater	carbohydrates
kollaps	collapse
kollapsade	collapsed
kollektiv	collective
kollektivtrafik	public
koloni	colony
koloniala	colonial
kolonialism	colonialism
kolonialismen	the colonialism
kolonialtiden	colonial
kolonier	colonies
kolonierna	colonies
kolonin	colony
koloniserades	colonized
koloniseringen	the colonization
kolväten	hydrocarbons
kom	came
koma	coma
kombattant	combatant
kombination	combination
kombinationen	combination
kombinationer	combinations
kombinerad	combined
kombinerade	combined
kombineras	combined
kombinerat	combined
kometer	comets
komiker	comedian
komintern	comintern
komma	come
kommande	upcoming
kommendör	commander
kommentar	comment
kommentarer	comments
kommenterade	commented
kommer	is
kommersiell	commercial
kommersiella	commercial
kommersiellt	commercial
kommissionen	commission
kommit	come
kommitté	committee
kommittén	committee
kommun	municipality
kommunal	municipal
kommunala	municipal
kommunen	municipality
kommuner	municipalities
kommunerna	municipalities
kommunicera	communicate
kommunicerar	communicates
kommunikation	communication
kommunikationer	communications
kommunism	communism
kommunismen	communism
kommunismens	communism
kommunister	communists
kommunisterna	communists
kommunistisk	communist
kommunistiska	communist
kommunistpartiet	the communist party
kommunistpartiets	communist party
komplett	complete
komplex	complex
komplexa	complex
komplext	complex
komplicerad	complicated
komplicerat	complicated
komplikationer	complications
komponenter	components
kompositör	composer
kompositörer	composers
kon	group
koncentration	concentration
koncentrationsläger	concentration camp
koncentrerad	concentrated
koncentrerade	concentrated
koncept	concept
konflikt	conflict
konflikten	conflict
konflikter	conflicts
kong	kong
kongo	congo
kongokinshasa	kong kinshasa
kongress	congress
kongressen	congress
kongresspartiet	congress
konkret	concrete
konkreta	concrete
konkurrens	competition
konkurrensen	competition
konkurrerande	competing
konkurs	bankruptcy
konsekvens	consequence
konsekvenser	consequences
konsekvenserna	impact
konsekvent	consistent
konsensus	consensus
konsert	concert
konserten	concert
konserter	concerts
konserterna	concerts
konserthus	concert hall
konservatism	conservatism
konservatismen	conservatism
konservativ	conservative
konservativa	conservative
konsolen	bracket
konspirationsteorier	conspiracy theories
konst	art
konstant	constant
konstantin	konstantin
konstantinopel	constantinople
konstaterade	found
konsten	art
konstitution	constitution
konstitutionell	constitutional
konstitutionella	constitutional
konstitutionen	constitution
konstnär	artist
konstnären	artist
konstnärer	artists
konstnärlig	artistic
konstnärliga	artistic
konstruerade	constructed
konstruktion	construction
konstverk	artwork
konsubstantiation	consubstantiation
konsul	consul
konsumtion	consumption
konsumtionen	consumption
kontakt	contact
kontaktade	contacted
kontakten	contact
kontakter	contacts
kontinent	continent
kontinentala	continental
kontinenten	continent
kontinentens	continent
kontinenter	continents
kontinuerlig	continuous
kontinuerligt	continuous
konto	account
kontor	office
kontrakt	contract
kontraktet	contract
kontrast	contrast
kontroll	control
kontrollen	control
kontrollera	control
kontrollerade	controlled
kontrollerar	controlling
kontrolleras	controlled
kontroverser	controversies
kontroversiell	controversial
kontroversiella	controversial
kontroversiellt	controversial
konung	king
konungarike	kingdom
konungariket	kingdom
konventionella	conventional
konventionen	convention
konventioner	conventions
konvertera	convert
konverterade	converted
kopia	copy
koppar	copper
koppla	connect
kopplad	connected to
kopplade	connected
kopplas	connected
kopplat	coupled; connected
koppling	coupling
kopplingar	connections
kopplingen	coupling
koprolali	coprolalia
koranen	the koran
korea	korea
koreakriget	the korean war
koreanska	korean
korn	grain
korrekt	correct
korrekta	correct
korruption	corruption
korruptionsindex	corruption index
kors	cross
korset	cross
kort	short
korta	short
kortare	shorter
kosmiska	cosmic
kosovo	kosovo
kosovos	kosovo
kostade	cost
kostar	costs
kostnaden	cost
kostnader	costs
kostnaderna	costs
kostym	costume
kr	kronas
kraft	force
kraften	force
krafter	forces
kraftfull	powerful
kraftig	strong
kraftiga	strong
kraftigare	stronger
kraftigt	heavily
kraftverk	power plant
krav	requirement
kraven	claims
kravet	claim
kreativitet	creativity
krets	circuit
kretsar	circles
kretsen	circuit
krig	war
krigare	warrior
krigen	wars
kriget	war
krigets	war
krigsmakt	armed forces
krigsmakten	armed forces
krigsslutet	war
kriminella	criminals
kring	around
kris	crisis
krisen	crisis
kriser	crises
kristen	christian
kristendom	christianity
kristendomen	christianity
kristendomens	christian
kristi	christ
kristian	kristian
kristiansson	kristiansen
kristinas	kristina's
kristna	christian
kristus	christ
krita	chalk
kriterier	criteria
kriterierna	criteria
kritik	criticism
kritiken	criticism
kritiker	critics
kritikerna	critics
kritiserade	criticized
kritiserades	criticized
kritiserar	criticize
kritiserat	criticized
kritiserats	criticized
kritisk	critical
kritiska	critical
kritiskt	critical
kroatien	croatia
kroatiens	croatian
kroatiska	croatian
kromosom	chromosome
kromosomer	chromosomes
kromosomerna	chromosomes
krona	crown
kronan	crown
kronisk	chronic
kroniska	chronic
kronor	kronor
kronprins	crown prince
kronprinsen	crown prince
kronprinsessan	crown princess
kropp	body
kroppar	bodies
kroppen	body
kroppens	body
krossa	crush
kryddor	spices
kräva	demand
krävde	required
krävdes	were required
kräver	requires
krävs	required
krävt	required
krönika	chronicle
kröntes	crowned
kub	cube
kuba	cuba
kubanska	cuban
kubas	cuba
kuben	cube
kuiperbältet	the kuiper belt
kulmen	the acme
kulminerade	culminated
kultur	culture
kulturarv	heritage
kulturell	cultural
kulturella	cultural
kulturellt	cultural
kulturen	culture
kulturer	cultures
kunde	could
kunder	customer
kung	king
kungafamiljen	royal family
kungahuset	royal family
kungamakten	monarchy
kungar	kings
kungariket	kingdom
kungarna	kings
kungen	king
kungens	king
kunglig	royal
kungliga	royal
kunna	to
kunnat	could
kunskap	knowledge
kunskapen	knowledge
kunskaper	knowledge
kupol	dome
kupp	coup
kurder	kurds
kurderna	kurds
kurdisk	kurdish
kurdiska	kurdish
kurdistan	kurdistan
kurfursten	elector
kuriosa	bric-a-brac
kurs	course
kurt	kurt
kusin	cousin
kust	coastal
kusten	coast
kuster	coasts
kusterna	coasts
kustlinje	coastline
kuwait	kuwait
kvadratkilometer	square kilometer
kvalificerade	qualifying
kvalitet	quality
kvar	left
kvarstod	remaining
kvarstår	remains
kvarter	block
kvarteret	block
kvartsfinalen	quarter finals
kvarvarande	remaining
kvast	broom
kvicksilver	quicksilver
kvinna	woman
kvinnan	woman
kvinnans	woman
kvinnlig	female
kvinnliga	female
kvinnor	women
kvinnorna	women
kvinnornas	women
kvinnors	women
kväll	evening
kvällen	hours
kväve	nitrogen
kyla	cold
kyrilliska	cyrillic
kyrka	church
kyrkan	church
kyrkans	church
kyrkliga	church
kyrkor	churches
kyrkorna	churches
kyros	cyrus
källa	source
källan	source
källkod	source code
källor	source
källorna	the sources
kämpa	fight
känd	known
kända	known
kände	felt
känna	feel
kännedom	knowledge
känner	know
kännetecken	characteristics
kännetecknas	characterized
känns	feels
känsla	feeling
känslan	sense
känslig	susceptible
känsliga	1st&2nd: fragile 3rd: sensitive
känslor	feelings
känt	known
kär	in love
kärlek	love
kärleken	the love
kärna	core
kärnan	core
kärnkraft	nuclear power
kärnkraftverk	nuclear power plant
kärnor	cores
kärnvapen	nuclear weapons
köket	cuisine
köln	köln
kön	sex
könen	the sexes
könsorgan	genitals
könsorganen	sex organs
köp	buy
köpa	buy
köpenhamn	copenhagen
köpenhamns	copenhagen
köper	buy
köpmän	merchants
köpt	purchased
köpte	bought
kör	drive
köra	drive
körberg	körberg
körs	run
kött	meat
l	l
la	la
laboratorium	laboratory
ladda	load
laddade	charged
laddning	charge
lade	added
lades	put
ladin	ladin
lag	law
lagar	laws
lagarna	laws
lagen	act
lager	stock
lagerkvist	lagerkvist
lagerlöf	lagerlöf
laget	team
lagets	side
lagförslag	bill
lagliga	legal
lagras	stored
lagring	storage
lagstiftande	legislative
lagstiftning	legislation
lagstiftningen	legislation
lagt	added
lagts	sent
laila	laila
lake	lake
land	country
landet	country
landets	its
landområden	land
lands	country
landsbygden	rural area
landshövding	governor
landskap	landscape
landskapen	provinces
landskapet	landscape
landskommun	rural municipality
landslag	national team
landslaget	football
landsting	county
lanka	lanka
lanserade	launched
lanserades	launched
lanseringen	release
laos	laos
larry	larry
lars	lars
larsson	larsson
larssons	larsson
laryngoskop	laryngoscope
lasse	lasse
lastbilar	trucks
lat	methacrylate
latin	latin
latinamerika	latin america
latinamerikanska	latin-american
latinet	latin
latinets	latin
latinska	latin
laura	laura
lava	lava
lawrence	lawrence
le	smile
led	point
leda	lead
ledamot	member
ledamöter	members
ledamöterna	members
ledande	leading
ledare	leader
ledaren	leader
ledarna	conductors
ledarskap	leadership
ledda	led
ledde	led
leddes	passed
leden	joint
leder	leads
ledger	ledger
ledning	management
ledningen	the lead
leds	passed
lee	lee
leeds	leeds
left|px	left px
legat	layed
legend	legend
legenden	legend
legender	legends
legitimitet	legitimacy
leipzig	leipzig
lejon	lion
lejonet	lion
lena	lena
lenin	lenin
lenins	lenin
lennart	lennart
lennon	lennon
leo	leo
leonard	leonard
leonardo	leonardo
leopold	leopold
les	les
let	let
leta	search
lett	resulted
lettland	latvia
leukemi	leukemia
lev	lev
leva	live
levande	live
levde	survived
lever	living
levern	the liver
levnadsstandard	standard of living
levnadsstandarden	living standard
levt	lived
lewis	lewis
lexikon	dictionary
liam	liam
libanon	lebanon
liberala	liberal
liberaler	liberals
liberalism	liberalism
liberalismen	liberalism
liberty	liberty
library	library
libyen	libya
lida	suffer
lidande	suffering
lider	suffer
lidit	suffered
liechtenstein	liechtenstein
life	life
liga	league
ligacupen	league cup
ligan	league
ligga	lie
liggande	lie
ligger	lies
light	light
lik	like
lika	equal
likartade	similar
likaså	also
likhet	similarity
likheter	similarities
liknade	similar
liknande	similar
liknar	similar
liknas	likened
liksom	as well as
likt	like
likväl	nevertheless
likör	liqueur
lilla	small
lima	lima
lina	line
lincoln	lincoln
linda	wind
lindgren	lindgren
lindgrens	lindgren
lindh	lindh
linje	line
linjen	line
linjer	lines
linjerna	lines
linköping	linköping
linköpings	linköping
linné	linneus
linux	linux
lisa	lisa
lisbet	lisbet
lissabon	lisbon
lissabonfördraget	lisbon treaty
list	cunning
lista	list
listade	listed
listan	list
listor	lists
listorna	menus
litauen	lithuania
lite	little
liten	small
liter	liters
litet	small
litteratur	literature
litteraturen	literature
litterär	literary
litterära	literary
liv	life
livealbum	live album
liverpool	liverpool
liverpools	liverpool
livet	life
livets	life
livslängd	life
livsmedel	food
livsstil	lifestyle
livstid	lifetime
liza	liza
ljud	sound
ljudet	sound
ljung	heather
ljungström	ljungström
ljus	light
ljusare	lighten
ljuset	light
locka	tempt
lockar	curls
locke	locke
loggbok	logbook
logik	logic
logotyp	logotype
lois	lois
lojalitet	loyality
lokal	local
lokala	local
lokaler	facilities
lokalt	local
london	london
londons	london
lopp	race
loppet	the race
lord	lord
loss	unstuck
lost	lost
lotta	lotta
louis	louis
louise	louise
louisiana	louisiana
lovade	promised
lovat	promised
lp	lp
lsd	lsd
lucas	lucas
lucia	lucia
lucky	lucky
ludvig	ludvig
ludwig	ludwig
luft	air
luften	air
lugn	quiet
lugna	calm
lukas	lukas
luleå	luleå
luminositet	luminosity
lundell	lundell
lundgren	lundgren
lunds	lund's
lunginflammation	pneumonia
lungorna	the lungs
lupus	lupus
lust	desire
luther	luther
luthers	luther
lutherska	lutheran
lutning	incline
luxemburg	luxemburg
lycka	happiness
lyckade	successful
lyckades	managed
lyckan	happiness
lyckas	succeed
lyckats	succeeded
lyder	obeys
lyfta	lift
lyfter	lifts
lyrik	poetry
lysande	brilliant
lyssna	listen
lyssnade	listened
lyssnar	listens
läge	location
lägenhet	apartment
läger	camp
läget	position
lägga	lay
läggas	added
lägger	put
läggs	added
lägre	lower
lägret	camp
lägst	lowest
lägsta	lowest
läkare	doctor
läkaren	doctor
läkemedel	drug
läkemedelsverket	medicines work
lämna	leave
lämnade	left
lämnades	left
lämnar	leaves
lämnas	left
lämnat	left
lämningar	remnants
lämplig	suitable
lämpliga	suitable
lämpligt	suitable
län	county
länder	countries
länderna	countries
ländernas	states
länders	countries
längd	length
längden	length
länge	long
längre	longer
längs	along
längst	farthest
längsta	longest
längtan	longing
länk	link
länkar	link
läns	county
lär	learn
lära	teach
läran	teaching
lärare	teacher
lärda	literate
lärde	learned
lärjungar	disciples
läror	teachings
lärt	learned
läs	read
läsa	read
läsare	reader
läsaren	reader
läser	reads
läses	read
läsning	reading
läst	read
läste	read
lät	made
lätt	easy
lätta	light
lättare	lighter
låg	low
låga	low
lågt	low
lån	loan
låna	borrow
lånat	borrowed
lång	long
långa	long
långbåge	long bow
långfilm	feature
långhårig	long-haired
långsamma	slow
långsammare	slowly
långsamt	slowly
långt	far
långtgående	far-reaching
långvarig	prolonged
långvariga	long-standing
långvarigt	long
låt	song
låta	sound
låtar	songs
låtarna	songs
låten	song
låter	sounds
låtit	chair
låtskrivare	song writers
löfte	promise
löften	promises
lön	salary
löner	salaries
lönneberga	lönneberga
löpande	current
löper	run
lördagen	saturday
lösa	solve
lösas	solved
löser	solves
lösning	solution
lösningar	solutions
lösningen	solution
lösningsmedel	solvent
löst	solved
löstes	dissolved
mabel	mabel
machu	machu
madagaskar	madagascar
madeira	madeira
madeleine	madeleine
madonna	madonna
madrid	madrid
maffia	mob
maffian	mob
magdalena	magdalena
magic	magic
magnetfält	magnetic field
magnetiska	magnetic
magnitud	magnitude
magnus	magnus
magnusson	magnusson
mahatma	mahatma
maiden	maiden
maidens	maidens
main	main
maj	may
majoritet	majority
majoriteten	majority
majs	corn
makadam	macadam
make	husband
makedonien	macedonia
makedonska	macedonian
makt	power
makten	power
maktens	forces
makter	powers
malaysia	malaysia
malcolm	malcolm
malin	malin
malmö	malmö
malmös	malmö
malta	malta
mamma	mother
man	man
manager	manager
manchester	manchester
mandat	mandate
mandatperiod	term
mandelas	mandelas
mando	command
manhattan	manhattan
mani	mania
maniska	manic
mankell	mankell
manlig	male
manliga	male
mannen	art
mannens	man
mans	male
manson	manson
manteln	the mantle
manuel	manuel
manus	script
manuskript	script
mao	mao
maos	maos
marco	marco
marcus	marcus
margaret	margaret
maria	maria
marie	marie
mariette	mariette
marijuana	marijuana
marilyn	marilyn
marina	marine
marinen	navy
marino	marino
mario	mario
marissa	marissa
mark	ground
markant	significant
marken	soil
markera	mark
markerade	selected
markerar	denotes
marklund	marklund
marknad	market
marknaden	market
marknader	markets
marknadsekonomi	market
markus	marcus
marley	marley
marleys	marley's
marocko	morocco
mars	march
marshall	marshall
martin	martin
marx	marx
marxism	marxism
marxismen	marxism
marxistisk	marxist
marxistiska	marxist
mary	mary
maskiner	machines
massa	mass
massachusetts	massachusetts
massakern	massacre
massan	mass
massiv	massive
massiva	massive
massmedia	mass media
massor	lots
master	master
mat	food
match	match
matchen	match
matcher	matches
matcherna	matches
matematik	mathematics
matematiken	mathematics
matematiker	mathematician
matematisk	mathematical
matematiska	mathematical
maten	the food
materia	matter
material	material
materialet	material
materiella	material
matrix	matrix
mats	mat's
matt	dull
matteus	matthew
matteusevangeliet	matthew
matthew	matthew
mattias	mattias
mattis	mattis
maurice	maurice
max	max
maya	maya
med	with
medan	while
medarbetare	coworker
medborgare	national
medborgarna	citizens
medborgarskap	citizenship
medborgerliga	civil
meddelade	announced
meddelande	message
meddelanden	messages
medel	average
medelhavet	mediterranean sea
medelhavsklimat	mediterranean climate
medelhavsområdet	the mediterranean region
medelklassen	middle class
medellivslängd	average lifespan
medeltemperaturen	the average temperature
medeltid	the medieval times
medeltida	medieval
medeltiden	middle ages
medeltidens	medieval
medelålder	middle age
medför	entails
medföra	result
medförde	resulted
medfört	resulted
media	media
medicin	medicine
mediciner	drugs
medicinering	medication
medicinsk	medical
medicinska	medical
medicinskt	medical
medier	media
mediet	medium
medina	medina
medlem	member
medlemmar	members
medlemmarna	members
medlemskap	membership
medlemsstat	member
medlemsstater	member
medlemsstaterna	member
medlemsstaternas	member
medverka	contribute
medverkade	participated; contributed
medverkan	participation
medverkar	involved
medverkat	participated
medvetande	consciousness
medveten	aware
medvetet	consciously
medvetna	conscious
mekaniska	mechanical
mekka	mecka
melankoli	melancholy
melker	melker
mellan	between
mellanfot	metatarsus
mellankrigstiden	interwar years
mellanrum	gap
mellanöstern	eastern
mellersta	middle
melodier	melodies
melodifestivalen	eurovision song contest
memoarer	memoirs
memorial	memorial
men	but
menade	meant
menar	mean
menas	means
menat	meant
mengele	mengele
mening	sentence
meningar	sentences
mental	mental
mentala	mental
mer	more
mera	more
mercurys	mercury
merkurius	mercury
merparten	most
merry	merry
mesopotamien	mesopotamia
messi	messi
messias	messiah
mest	most
mesta	most
mestadels	mostly
metabolism	metabolism
metaforer	metaphors
metall	metal
metaller	metals
metallica	metallica
metan	methane
meter	meter
metionin	methionine
metod	method
metoden	method
metoder	methods
metro	metro
mexico	mexico
mexikanska	mexican
mexiko	mexico
meyer	meyer
mfl	etc
miami	miami
michael	michael
michail	michail
michel	michel
michelle	michelle
michigan	michigan
mick	mike (microphone)
microsoft	microsoft
midsommar	midsummer
mig	me
miguel	miguel
mikael	mikael
mike	mike
mil	mil
milan	milan
milano	milano
mild	mild
milda	mild
mildare	milder
miley	miley
militär	military
militära	military
militären	military
militärer	soldiers
militärt	military
miljard	billion
miljarder	billions
miljon	million
miljoner	million
miljontals	millions
miljö	environment
miljöer	environments
miljön	the environment
miljöproblem	environmental problems
miller	miller
milt	mild
min	my
mina	mine
mind	mind
mindre	less
mineral	mineral
mineraler	minerals
miniatyr	miniature
miniatyr|	miniature
miniatyr|en	thumbnail
miniatyr|karta	thumbnail map
miniatyr|px|den	miniature
miniatyr|px|en	miniature
miniatyr|px|ett	miniature
minister	minister
ministerrådet	ministers
ministrar	ministers
minne	memory
minnen	memories
minnet	memory
minns	remember
minoritet	minority
minoriteten	minority
minoriteter	minorities
minoritetsspråk	minority
minska	reduce
minskad	reduced
minskade	decreased
minskar	decrease
minskat	reduced
minskning	reduction
minst	at least
minsta	minimum
minut	minute
minuter	minutes
miss	miss
missbruk	abuse
missförstånd	misunderstanding
misshandel	assault
mission	mission
missionärer	missions
misslyckade	failed
misslyckades	failed
misslyckande	failure
misslyckas	fail
misslyckats	failed
missnöje	dissatisfaction
missnöjet	discontent
misstag	mistake
misstänkt	suspected
misstänkta	suspected
mitt	my
mitten	middle
mix	mix
mjölk	milk
mm	millimeter
moberg	moberg
mod	courage
mode	fashion
modell	model
modellen	model
modeller	models
moder	mother
moderata	moderate
moderaterna	moderates
modern	modern
moderna	modern
modernare	more modern
modernismen	modernism
modernistiska	modernistic
modernt	modern
modersmål	mother tongue
modet	courage
modo	modo
mohammed	mohammed
moldavien	moldova
molekyler	molecules
moln	cloud
mona	mona
monaco	monaco
monark	monarch
monarken	monarch
monarki	monarchy
monarkin	monarchy
monetära	monetary
mongoliet	mongolia
monica	monica
monicas	monica
monografi	monograph
monopol	monopoly
monoteism	monotheism
monoteistiska	monotheistic
monroe	monroe
monster	monster
montana	montana
monte	assembly
montenegro	montenegro
monument	monument
moore	moore
mor	mother
mora	mora
moral	morality
moralisk	moral
moraliska	moral
moraliskt	morally
mord	murder
morden	murder
mordet	murder
morgan	morgan
morgon	morning
morgonen	morning
morris	morris
moseboken	genesis
moses	moses
moskva	moscow
mot	against
motion	exercise
motiv	subjects
motiveringen	the motivation
motivet	subject
motor	engine
motors	engine's
motorväg	motorway
motorvägar	highways
motorvägarna	the highways
motorvägen	motorway
motsats	contrast
motsatsen	the opposite
motsatt	opposite
motsatta	opposite
motsatte	opposed
motstånd	resistance
motståndare	opponents
motståndaren	the opponent
motståndarna	opponents
motståndet	the resistance
motståndsrörelsen	resistance
motsvarande	corresponding
motsvarar	corresponds
motsvarighet	equivalent
motsättningar	oppositions
mottagande	host
mottagare	receiver
mottagaren	receiver
mottagarens	receiver
motto	motto
mottog	received
motverka	counteract
mountain	mountain
movie	movie
mozart	mozart
mozarts	mozart
moçambique	mozambique
mr	mr
ms	motor ship
mtv	mtv
muhammad	muhammad
muhammed	muhammed
muhammeds	mohammed
mullusfiskar	goatfish
mun	mouth
munnen	mouth
mur	wall
muren	wall
murray	murray
muse	muse
museer	museums
museet	museum
museum	museum
music	music
musik	music
musikalen	musical
musikalisk	musical
musikaliska	musical
musikaliskt	musically
musiken	music
musikens	music
musiker	musicians
musikstil	music still
musikstilar	genres
musikvideo	music video
musikvideon	music video
musikvideor	music videos
muskler	muscles
musklerna	muscles
muslim	muslim
muslimer	muslims
muslimerna	muslims
muslimsk	muslim
muslimska	muslim
mussolini	mussolini
mussolinis	mussolini
mutationer	mutations
mycket	very
myndighet	authority
myndigheten	authority
myndigheter	authorities
myndigheterna	authorities
mynnar	opening
mynning	mouth
mynt	coin
myntade	coined
myntades	was coined
mysterium	mystery
mystiska	mystical
myter	myths
mytologi	mythology
mytologin	mythology
mytologiska	mythological
mäktiga	powerful
mäktigaste	most powerful
mälaren	mälaren
män	men
mängd	amount
mängden	amount
mängder	amounts
männen	men
människa	person
människan	the human
människans	human
människas	human
människor	people
människorna	people
människors	human
mänsklig	human
mänskliga	human
mänskligheten	humanity
mänsklighetens	human
mänskligt	human
märke	make
märken	brands
märks	labeled
märktes	labeled
märta	pain
mästare	master
mästarna	the champions
mäta	measure
mäter	measure
mätningar	measurements
mäts	measured
mätt	measured
må	feel
mål	case
måla	paint
målade	painted
målare	painter
målen	cases
måleri	painting
målet	the target
målning	painting
målningar	paintings
målningen	milling
målvakt	goalkeeper
målvakten	goalkeeper
mån	concerned
månad	month
månaden	month
månader	months
månaderna	months
månar	moons
månarna	moons
måne	moon
månen	moon
månens	the moon's
många	many
mångfald	diversity
måste	must
mått	measure
möjlig	possible
möjliga	possible
möjligen	possibly
möjliggjorde	made possible
möjliggör	enables
möjlighet	ability
möjligheten	the possibility
möjligheterna	possibilities
möjligt	possible
mönster	pattern
mördad	murdered
mördade	killed
mördades	killed
mörk	dark
mörkare	darker
mörker	darkness
mörkt	dark
möta	meet
möte	meeting
möten	meetings
möter	face
mötet	meeting
mötley	mötley
möts	met
mött	met
mötte	met
möttes	met
münchen	munich
n	n
nacka	nacka
nagasaki	nagasaki
namibia	namibia
namn	name
namnen	names
namnet	the name
nancy	nancy
napoleon	napoleon
napoleons	napoleon
narkotika	drug
nasa	nasa
nash	nash
nathan	nathan
nation	nation
national	national
nationalencyklopedin	the national encyclopedia
nationalförsamlingen	national assembly
nationalism	nationalism
nationalismen	nationalism
nationalister	nationalists
nationalistiska	nationalistic
nationalitet	nationality
nationalpark	national park
nationalparker	national parks
nationell	national
nationella	national
nationellt	nationally
nationen	nation
nationens	nation
nationer	nations
nationerna	nations
nationernas	nations
nations	nation
nato	nato
natt	night
natten	overnight
nattetid	overnight
natur	nature
natural	natural
naturen	nature
naturens	nature
naturgas	natural gas
naturlig	natural
naturliga	natural
naturligt	natural
naturligtvis	course
naturresurser	natural resources
naturtillgångar	natural resources
naturvetenskapliga	science
nazismen	nazi
nazisterna	nazis
nazisternas	nazi
nazistiska	nazi
nazityskland	nazi germany
nazitysklands	nazi germany
ned	down
nedan	below
nederbörd	precipitation
nederbörden	precipitation
nederlag	defeat
nederländerna	netherlands
nederländska	dutch
nedgång	decline
nedre	lower
nedsatt	reduced
nedåt	down
need	need
negativ	negative
negativa	negative
negativt	negative
neil	neil
nej	no
nelson	nelson
neo	neo
neologi	neology
nepal	nepal
neptunus	neptune
ner	down
nere	down
nervosa	nervosa
nervsystemet	nervous system
neutral	neutral
neutrala	neutral
neutralitet	neutral
neutralt	neutral
neutroner	neutrons
nevada	nevada
newport	newport
newton	newton
newtons	newton
nf	nf
nhl	nhl
ni	you
nickel	nickel
nicklas	nicklas
niclas	niclas
nietzsche	nietzsche
nietzsches	nietzsche
nigeria	nigeria
nikki	nikki
niklas	niklas
nikola	nikola
nikolaj	nikolaj
nils	nils
nilsson	nilsson
nio	nine
nionde	ninth
nirvana	nirvana
nivå	level
nivåer	levels
nivån	level
nixon	nixon
njurarna	the kidneys
nku	nku
nobel	nobel
nobelkommittén	the nobel commitee
nobelpriset	the nobel prize
nobelpristagare	nobel laureate (-s); nobel prize winner (-s)
nobels	nobel
nobelstiftelsen	nobel foundation
nog	probably
noga	carefully
noll	zero
nominerad	nominated
nominerades	nominated
nomineringar	nominations
nord	north
nordafrika	north africa
nordamerika	north america
nordamerikanska	north american
norden	north
nordens	nordic
nordirland	north ireland
nordisk	nordic
nordiska	nordic
nordiskt	nordic
nordkorea	north korea
nordkoreanska	north korean
nordkoreas	north korea
nordliga	northern
nordligaste	northernmost
nordost	northeast
nordsjön	north sea
nordväst	northwest
nordvästra	northwest
nordöst	northeast
nordöstra	northeast
norge	norway
norges	norway
normal	normal
normala	normal
normalt	normally
norman	norman
normer	standards
norr	north
norra	north
norrköping	norrköping
norrköpings	norrköping
norrland	northern
norrlands	norrland
norrmän	norwegian
norrut	north
norsk	norwegian
norska	norwegian
norstedt	norstedt
norstedts	collins
north	north
notation	notation
noter	notes
notera	note
noterade	note
nou	nou
nova	nova
november	november
now	now
nr	no
nsdap	nsdap
nu	now
nuförtiden	nowadays
nukleotider	nucleotides
numera	nowadays
nummer	number
nutid	present
nutida	contemporary
nuvarande	current
ny	new
nya	new
nyare	newer
nybildade	newly formed
nye	new
nyfödda	newborn
nyheten	news
nyheter	news
nyligen	recently
nytt	new
nytta	benefit
nyval	new election
nämligen	namely
nämnas	mentioned
nämnda	said
nämnde	mentioned
nämner	mentions
nämns	mentioned
nämnts	mentioned
när	when
nära	near
närhet	closeness
näring	nutrition
näringsliv	business
näringslivet	business
närliggande	nearby
närma	approach
närmade	approached
närmar	close in
närmare	close to
närmast	closest
närmaste	closest
närstående	related
närvarande	present
närvaro	presence
näsan	the nose
näst	second
nästa	next
nästan	almost
nät	web
nätet	net
nätverk	network
nätvingar	neuroptera
nå	reach
nåd	grace
nådde	reached
nåddes	reached
någon	someone
någonsin	ever
någonstans	somewhere
någonting	anything
någorlunda	fairly
något	something
några	a few
når	reaches
nås	reached
nått	reached
nöd	need
nödvändig	necessary
nödvändiga	necessary
nödvändigt	necessary
nödvändigtvis	necessarily
nöjd	content
o	o
oavgjort	tie
oavsett	regardless
obama	obama
obamas	obama
obelix	obelix
oberoende	independent
objekt	object
objekten	items
objektet	object
obligatorisk	obligatory
obligatoriskt	mandatory
observationer	observations
observatörer	observers
observera	note
observeras	observed
oc	oc
oceanen	ocean
och	and
ocheller	and/or
också	also
ockupation	occupation
ockupationen	occupation
ockuperade	occupied
ockuperades	occupied
ockuperat	occupied
oden	oden
odens	odin's
odlade	cultured
odlas	cultured
odling	culture
oecd	oecd
oerhörd	enormous
oerhört	tremendously
of	of
off	off
offensiven	offensive
offentlig	public
offentliga	public
offentligt	publicly
offer	victims
office	office
officerare	officers
official	official
officiell	official
officiella	official
officiellt	officially
offren	victims
offret	victim
offside	offside
ofta	often
oftare	more often
oftast	usually
oförmåga	inability
ogillade	dismissed
oklart	clear
oktober	october
oktoberrevolutionen	october revolution
okänd	unknown
okända	unknown
okänt	unknown
ola	ola
olagligt	illegal
olika	different
oliver	olives
olja	oil
olle	olle
ollonet	glans
olof	olof
olsson	olsson
olycka	accident
olyckan	accident
olyckor	accidents
olympia	olympia
olympiastadion	olympa stadium
olympiska	olympic
om	if
ombord	onboard
omedelbar	immediate
omedelbart	immediately
omfatta	include
omfattade	included
omfattande	large
omfattar	encompass
omfattas	covered
omfattning	extent
omger	surrounds
omges	surrounded
omgivande	ambient
omgiven	surrounded
omgivning	environment
omgivningen	surroundings
omgående	immediately
omgångar	in turns; periods; mandates
omgången	round
omkom	died
omkring	about
omkringliggande	surrounding
omloppsbana	orbit
omloppsbanor	orbit
omnämns	mentioned
område	area
områden	area
områdena	regions
området	area
områdets	area
omröstning	vote
omröstningen	vote
omskärelse	circumcision
omslaget	cover
omstritt	controversial
omständigheter	circumstances
omtvistat	contentious
omvandlar	transmuted
omvandlas	converted
omvandling	conversion
omvända	reverse
omvänt	reversed
omvärlden	abroad
omväxlande	varied
omöjligt	impossible
on	on
onani	masturbation
onda	evil
ondska	evil
ondskan	evil
ont	evil
ontario	ontario
open	open
opera	opera
operan	opera
operation	operation
operationer	operations
operativsystem	os
opinion	opinion
opinionen	opinion
opposition	opposition
oppositionen	opposition
oralsex	oral sex
orange	orange
ord	words
ordagrant	literally
ordbok	dictionary
orden	words
ordentligt	proper
ordet	the word
ordförande	president
ordinarie	ordinary
ordna	arrange
ordnade	arranged
ordnar	fix
ordning	order
ordningen	the order
ordspråk	proverb
organ	organ
organisation	body
organisationen	organization
organisationens	organization
organisationer	organizations
organisera	organize
organiserad	organized
organiserade	organized
organiseras	organized
organiserat	organized
organisk	organic
organiska	organic
organism	organism
organismen	organism
organismer	organisms
orgasm	orgasm
origin	original
original	original
orkester	orchestra
ormar	snakes
oro	concern
orolig	worried
oroligheter	unrest
orsak	cause
orsaka	cause
orsakad	caused
orsakade	caused
orsakar	cause
orsakas	caused
orsakat	caused
orsaken	cause
orsaker	causes
orsakerna	causes
ort	city
orten	the suburb
orter	visited
ortodoxa	orthodox
os	os
oscar	oscar
oskar	oskar
oslo	oslo
osmanerna	ottoman turks
osmanska	osmanian
oss	center
ost	cheese
osv	etc
osäker	uncertain
osäkert	uncertain
osäkra	insecure
otaliga	countless
otto	otto
out	out
ovan	above
ovanför	above
ovanlig	unusual
ovanliga	rare
ovanligt	unusual
ovanpå	top
ovanstående	above
oväntat	unexpectedly
own	own
oxenstierna	the oxenstierna
oxford	oxford
ozzy	ozzy
oändligt	infinitely
pablo	pablo
page	page
pakistan	pakistan
palats	palace
palestina	palestine
palestinier	palestinian
palestinsk	palestinian
palestinska	palestine
palme	palme
palmes	palme's
pamela	pamela
panthera	panthera
pappa	dad
papper	paper
par	pair
paradiset	paradise
paraguay	paraguay
parallella	parallel
parallellt	parallel
parentes	brackets
paret	pair
paris	paris
park	park
parken	park
parker	parks
parlament	parliament
parlamentarisk	parliamentary
parlamentariska	parliamentary
parlamenten	parliaments
parlamentet	house
parlamentets	parliament
parlamentsvalet	parliamentary
parten	party
parter	parties
parterna	parties
parti	party
partido	partido
partier	portions
partierna	portions
partiet	party
partiets	party
partiklar	particles
partiledare	party leader
partner	partner
partnern	partner
pass	pass
passa	fit
passade	free
passagerare	passenger
passagerarna	passengers
passande	suitable
passar	suits
passera	pass
passerade	passed
passerar	pass
passiv	passive
pastor	pastor
pastoral	pastoral
patent	patent
patienten	the patient
patienter	patients
patrick	patrick
patrik	patrik
patterson	patterson
paul	paul
paulo	paulo
paulus	paul
paus	pause
paz	paz
pc	pc
peang	forceps
pearl	pearl
peka	point
pekar	point
pekat	identified
peking	beijing
pelle	pellet
pendeltåg	commuter
pengar	money
pengarna	the money
penis	penis
pennsylvania	pennsylvania
people	people
per	per
perfekt	perfect
performance	performance
period	period
perioden	period
perioder	period
periodiska	periodic
periodvis	periodically
permanent	permanent
permanenta	permanent
pernilla	pernilla
perro	perro
perry	perry
persbrandt	persbrandt
perserna	persian
persien	persian
persiska	persian
person	person
personal	staff
personalen	the staff
personen	person
personens	person
personer	people
personerna	people
personlig	personal
personliga	personal
personligen	personally
personlighet	personality
personlighetsstörning	personality
personlighetsstörningar	personality disorders
personligt	personally
persons	person
perspektiv	perspective
persson	persson
peru	peru
peruanska	peruvian
pest	plague
pesten	plague
peter	peter
peters	peters
petersburg	petersburg
petra	petra
petroleum	petroleum
petrus	peter
petter	petter
pettersson	pettersson
pga	"because of (short of ""på grund av"")"
ph	ph
phil	phil
philadelphia	philadelphia
philip	philip
philips	philips
phoebe	phoebe
phoenix	phoenix
pi	pi
piano	piano
picasso	picasso
picchu	picchu
picture	picture
pierre	pierre
pilatus	pilate
pink	pink
pippi	pippi
pippin	pippin
pirate	pirate
piratpartiet	pirate party
pitt	pitt
pjäs	play
pjäsen	piece
pjäser	plays
place	place
placera	place
placerad	placed
placerade	placed
placerades	placed
placerar	place
placeras	placed
placering	placement
plan	plan
planen	pitch
planer	plans
planerad	planned
planerade	planned
planerar	plans
planeras	planned
planerat	planned
planering	planning
planerna	plans
planet	planet
planeten	planet
planetens	planet
planeter	planets
planeterna	planets
planeternas	planets
plasma	plasma
platina	platinum
platon	platon
platons	platos
plats	place
platsen	place
platser	places
platt	flat
platta	plate
plattan	plate
plattform	platform
platån	plateau
player	player
playstation	playstation
plikt	duty
plikter	duties
plocka	pick
plural	plural
plus	plus
pluto	pluto
plötsligt	suddenly
poe	poe
poes	poe
poesi	poetry
poet	poet
poeten	poet
poeter	poets
point	point
pojkar	boys
pojkarna	boys
pojke	boy
pojkvän	boyfriend
polacker	poles
polen	poland
polens	polands
policy	policy
polis	police
polisen	police
polisens	police
poliser	police
politik	policy
politiken	policy
politiker	politician
politisk	political
politiska	political
politiskt	political
polska	polish
pommern	pommern
pompejus	pompejus
ponny	pony
pontus	pontus
pop	pop
popsångare	pop singer
popularitet	popularity
population	population
populationen	population
populationer	populations
populär	popular
populära	popular
populäraste	nearby
populärkultur	popular
populärkulturen	popular culture
populärmusik	popular
populärt	popularly
port	port
porto	postage
porträtt	portrait
portugal	portugal
portugals	portugals
portugisiska	portuguese
position	position
positionen	position
positioner	positions
positiv	positive
positiva	positive
positivt	positive
post	not a swedish word
posten	the position
poster	items
postumt	posthumously
potatis	potato
potential	potential
potentiellt	potential
potter	potter
povel	povel
poäng	point
prag	prague
praktiken	practice
praktisk	practical
praktiska	practical
praktiskt	practically
prata	talk
pratar	talking
praxis	practice
precis	just
premier	premiums
premiär	premiere
premiären	premiere
premiärminister	prime minister
premiärministern	the prime minister
preparat	substance
presenterade	presented
presenterades	presented
presenterar	presents
presenteras	presented
president	president
presidenten	president
presidentens	the president's
presidenter	presidents
presidentvalet	presidential elections
presley	presley
press	press
pressas	pressed
pressen	press
prestigefyllda	prestigious
preussen	prussia
preventivmedel	contraceptives
primitiva	primitive
primtal	prime number
primära	primary
prince	prince
princip	principle
principen	principle
principer	principles
prins	prince
prinsen	prince
prinsessan	princess
pris	award
priser	prices
priserna	prices
priset	price
prisma	prism
pristagare	laureate
privat	private
privata	private
privatliv	private
privilegier	privileges
privilegium	privilege
problem	problem
problemen	problems
problemet	the problem
procent	percent
process	process
processen	process
processer	processes
producent	producer
producenten	producer
producenter	producers
producera	produce
producerad	produced
producerade	produced
producerades	produced
producerar	producing
produceras	produced
producerat	produced
producerats	produced
produkt	product
produkten	product
produkter	products
produktion	production
produktionen	production
produktiv	productive
professionell	professional
professionella	professional
professor	professor
professorn	professor
profet	prophet
profeten	prophet
profeter	prophet
profil	profile
programledare	host
programmet	the program
programvara	software
projekt	project
projektet	project
prokaryoter	prokaryote
promemoria	memorandum
propaganda	propaganda
proportioner	proportions
prosa	prose
protein	protein
proteiner	proteins
proteinerna	proteins
proteinet	protein
protestanter	protestants
protestantiska	protestant
protester	protests
protesterade	protested
protesterna	protests
protokoll	protocol
protoner	protons
prov	tests
provins	province
provinsen	province
provinser	provinces
provinserna	provinces
provisoriska	provisional
prägel	character
präglad	characterized
präglade	characterized
präglades	was marked
präglas	characterized
präglats	characterized
präster	priests
ps	ps
psykisk	psychological
psykiska	psychic
psykiskt	psychic
psykologi	psychology
psykologin	psychology
psykologisk	psychological
psykologiska	psychological
psykos	psychosis
psykosen	psychosis
psykoser	psychoses
psykoterapi	psychotherapy
psykotiska	psychotic
publicera	publish
publicerad	published
publicerade	published
publicerades	published
publiceras	published
publicerat	published
publiceringen	publishing
publik	audience
pucken	the puck
puerto	puerto
puls	pulse
pund	pound
punk	punk
punkt	point
punkten	point
punkter	points
purple	purple
pythagoras	pythagoras
päls	fur
pär	pär
på	on
påbörjade	started
påbörjades	started
påbörjas	starts
påföljande	subsequent
pågick	went
pågående	ongoing
pågår	(in) progress
påminde	reminded
påminner	reminds
påsk	easter
påsken	easter
påstod	claimed
påstådda	alleged
påstående	statement
påståenden	claims
påstår	states
påstås	claimed
påtagligt	substantially
påtryckningar	pressure
påven	the pope
påverka	affect
påverkad	affected
påverkade	affected
påverkades	affected
påverkan	impact
påverkar	affect
påverkas	affected
påverkat	affected
påverkats	affected
påvisa	prove
q	q
queen	queen
queens	queen
rachel	rachel
rachels	rachel
rad	row
radie	radius
radikala	radical
radikalt	radically
radio	radio
radioaktiva	radioactive
radioaktivt	radioactive
radion	radio
rafael	rafel
ragnar	ragnar
raid	raid
rainbow	rainbow
rak	straight
raka	straight
rakt	straight
ramadan	ramadan
ramel	frame
ramels	ramel's
ramen	frame
rammstein	rammstein
rankas	ranks
rankning	ranking
rankningar	rankings
rapport	report
rapporten	report
rapporter	reports
rapporterade	reported
rapporterar	reports
ras	race
rasade	collapsed
rasen	breed
raser	species
rasism	racism
rastafari	rastafarian
rastafarianer	rastafarian
rastafarianerna	the rastafarian
reagan	reagan
reagans	reagan
reagera	reacting
reagerar	reacts
reaktion	reaction
reaktionen	reaction
reaktioner	reactions
reaktionerna	reactions
reaktorer	reactors
reaktorn	reactor
realiteten	positive
rebecca	rebecca
recensioner	reviews
receptorer	receptors
red	ed
reda	find out
redaktör	editor
redan	already
rede	nest
rederiet	the shipping company
redo	ready
redovisas	reported
redskap	gear
reducera	reduce
reduktion	reduction
referens	reference
referenser	references
refererar	refers
reform	reform
reformationen	the reformation
reformer	reforms
regel	rule
regelbunden	regular
regelbundet	regularly
regelbundna	regular
regeln	rule
regent	regent
regenter	monarchs
regerade	ruled
regerande	ruling
regering	government
regeringar	governments
regeringen	government
regeringens	government
regeringschef	government
regeringsmakten	the government
regeringstid	term of government
reggae	reggae
reggaen	reggae
regi	direction
regim	regime
regimen	regime
regimer	regimes
region	region
regional	regional
regionala	regional
regionalt	regional
regionen	region
regioner	regions
regionerna	regions
regisserad	directed
regissör	director
regissören	director
registrerade	recorded
regler	regulations
reglera	controlling
reglerar	regulates
regleras	controlled
reglerna	rules
regn	rain
regnar	rain
regnskog	rainforest
reguljära	regular
reidar	reidar
reidars	reidars
reinfeldt	reinfeldt
reklam	advertising
reklamen	ad
rekord	record
rekordet	record
relaterade	related
relation	relationship
relationen	relationship
relationer	relationships
relationerna	relations
relativa	relative
relativt	relatively
releasedatum	released
religion	religion
religionen	religion
religionens	religion
religioner	religions
religionerna	religions
religionsfrihet	religion
religiös	religious
religiösa	religious
religiöst	religious
remmer	remmer
ren	clean
rena	clean
rent	true
renässans	renaissance
renässansen	renaissance
rené	rené
reologi	rheology
reportrar	reporters
representant	representative
representanter	representatives
representanthuset	representatives
representation	representation
representativ	representative
representera	represent
representerade	represented
representerar	represents
representeras	represented
reptiler	reptiles
republik	republic
republika	republic
republikanska	republican
republiken	republic
republikens	republic
republiker	republics
resa	travel
resan	the trip
resande	travelling
research	research
reser	travels
residensstad	county
resolution	resolution
resor	travels
respekt	respect
respektive	respective
rest	remain
restaurang	restaurant
restauranger	restaurants
reste	traveled
resten	rest
rester	remains
resterande	remaining
resultat	results
resultaten	results
resultatet	result
resultera	result
resulterade	resulted
resulterar	results
resulterat	resulted
resurs	resource
resurser	resources
retorik	rhetoric
retoriken	rhetoric
retoriska	rhetorical
revir	territory
revolution	revolution
revolutionen	revolution
revolutionens	revolution
revolutionär	revolutionary
revolutionära	revolutionary
revs	was demolished
reza	reza
rhen	the rhine
rice	rice
richard	richard
richards	richards
richmond	richmond
rico	rico
riddare	knight
rik	rich
rika	rich
rikare	richer
rikaste	richest
rike	kingdom
rikedom	wealth
riken	kingdoms
riket	kingdom
rikets	its
riksdag	parliament
riksdagen	parliament
riksdagens	parliament
riksdagsvalet	parliament election
riksförbundet	national association
rikskansler	chancellor
riksrådet	privy council; council of state; crown council; senate
riksväg	highway
rikt	rich
riktad	directed
riktade	directed
riktar	target
riktas	directed
riktat	directed
riktig	true
riktiga	real
riktigt	really
riktlinjer	guidelines
riktning	direction
riktningar	directions
riktningen	direction
ring	ring
ringa	call
ringar	rings
ringde	called
ringen	ring
rinner	flows
ris	rice
risk	risk
risken	the risk
risker	risks
riskerar	risk
rita	draw
ritualer	rituals
rivalitet	rivalry
river	river
rna	rna
rob	rob
robbie	robbie
robert	robert
roberto	roberto
roberts	roberts
robin	robin
robinson	robinson
rockband	rock band
rocken	the rock
rockgrupper	rock groups
rocksångare	rock singer
rod	rod
roger	roger
roland	roland
roll	role
rollen	role
roller	roles
rollfigur	character
rollfigurer	characters
rolling	rolling
rom	rome
roma	roma
roman	novel
romance	romance
romanen	novel
romaner	novels
romani	romani
romantiken	romance
romantikens	romantic
romantiska	romantic
romarna	the roman
romarriket	the roman empire
romeo	romeo
romer	romani people
romerna	roma
romersk	roman
romerska	roman
romerske	roman
romerskkatolska	roman catholic
roms	rome's
romska	romani
romulus	romulus
ron	rose
ronaldinho	ronaldinho
ronaldo	ronaldo
ronden	round
ronja	ronja
roosevelt	roosevelt
rorsman	helmsman
rosa	pink
rose	rose
rosenberg	rosenberg
rotation	rotation
roterande	rotating
roterar	rotates
rousseau	rousseau
rovdjur	predator
rowling	rowling
roy	roy
rubiks	rubik's
rubrik	heading
rudolf	rudolf
rugby	rugby
ruiner	ruins
rum	room
rummet	room
rumänien	romania
rumänska	romanian
run	run
runda	round
running	running
runor	runes
runorna	runes
runstenar	runestones
runt	around
runtom	around
ruset	the fuddle
rush	rush
russell	russell
rwanda	rwanda
ryan	ryan
rybak	rybak
rygg	back
ryggen	back
rykte	reputation
rykten	rumors
rymden	space
rymmer	hold
rysk	russian
ryska	russian
ryssland	russia
rysslands	russian
rytmiska	rhythmic
räcker	enough
räckte	handed
rädd	afraid
rädda	save
räddade	saved
räddar	saves
rädsla	fear
räkna	count
räknade	calculated
räknar	counts
räknas	calculated
räknat	calculated
rätt	right
rätta	correct
rättegång	trial
rättegången	trial
rätten	right
rätter	dishes
rättigheter	rights
rättigheterna	rights
rättsliga	legal
rättvisa	justice
råd	advice
rådande	current
rådde	prevailed
råder	is
rådet	the council
rådets	council
rådgivare	advisor
rådhus	town hall
råkar	happens to
råolja	crude oil
råvaror	raw
röd	red
röda	red
röka	smoke
rökning	smoking
rör	touch, move(-s)
röra	move
rörande	concerning
rörde	touched
rörelse	movement
rörelsen	movement
rörelsens	movement
rörelser	movements
rörelserna	the movements
rörlighet	movement
röst	voice
rösta	vote
röstade	voted
rösten	voice
röster	votes
rösterna	votes
rösträtt	vote
rött	red
rötter	roots
sa	said
saab	saab
sabbath	sabbath
sachsen	saxony
saddam	saddam
sade	said
sades	said
saga	saga
sagan	tale
sagor	tales
sagt	said
sahara	sahara
sahlin	sahlin
saint	saint
sak	thing
saken	matter
saker	things
saknade	missing
saknades	missing
saknar	lacks
saknas	missing
sakrament	sacrament
sakta	slowly
salt	salt
salvador	salvador
sam	co
samarbeta	cooperate
samarbetade	collaborated
samarbetar	collaborates
samarbetat	collaborated
samarbete	cooperation
samarbeten	co
samarbetet	co
samband	connection
sambandet	connection
same	same
samerna	the lapp
samfund	society
samfundet	community
samhälle	society
samhällen	communities
samhället	society
samhällets	society
samisk	sami
samiska	sami
samla	collect
samlade	collected
samlades	gathered
samlag	intercourse
samlar	collect
samlat	collected
samlats	collected
samling	collection
samlingar	collections
samlingsalbum	compilations
samma	same
samman	together
sammanfaller	coincides
sammanfattning	summary
sammanhang	context
sammanhanget	context
sammanhängande	continous
sammanlagt	total
sammansatt	composed
sammansatta	composed
sammansättning	composition
samoa	samoa
samspel	interaction
samt	and
samtal	call
samtida	contemporary
samtidigt	while
samtliga	all
samtycke	approval
samuel	samuel
samverkan	cooperation
samverkar	co
samväldet	commonwealth
san	san
sand	sand
sandy	sandy
sankt	sankt
sankta	saint
sann	true
sanna	true
sanning	truth
sanningen	truth
sannolikhet	probability
sannolikt	likely
sanskrit	sanskrit
sant	true
santa	santa
santiago	santiago
sapiens	sapiens
sara	sara
sarah	sarah
sarajevo	sarajevo
satan	devil
satanism	satanism
sats	clause
satsa	bet
satsade	bet
satsningar	investments
satt	sat
satte	sat
sattes	added
saturnus	saturnus
saudiarabien	saudi arabia
sauron	sauron
sawyer	sawyer
scen	scene
scenen	stage
scener	scenes
schack	chess
schizofreni	schizophrenia
schwarzenegger	schwarzenegger
schweiz	switzerland
schweiziska	swiss
science	fiction
scientologikyrkan	the church of scientology
scott	scott
screen	screened
se	see
sean	sean
sebastian	sebastian
sed	custom
sedan	then
sedd	seen
seden	custom
seder	subsequently
sedermera	subsequently
sedlar	bills
seger	win
segern	win
seglade	sailed
segrar	wins
sekel	century
sekelskiftet	turn
sekreterare	secretary
sekt	sect
sekter	sects
sektion	section
sektorn	sector
sekulär	secular
sekulära	secular
sekunder	seconds
sekvens	sequence
selassie	selassie
selma	selma
semifinal	semi finals
semifinalen	semi finals
sen	late
sena	late
senare	later
senast	last
senaste	last
senaten	senate
senator	senator
sent	late
sentida	recent
separat	separate
separata	separate
separerade	separated
september	september
ser	see
serber	serbs
serbien	serbia
serbiens	serbia
serbisk	serbian
serbiska	serbian
serie	series
serien	series
seriens	series
serier	series
serotonin	serotonin
serveras	is served
service	service
servrar	servers
ses	be
seth	seth
sett	seen
setts	observed
sevärdheter	attractions
sex	six
sexton	sixteen
sexualitet	sexuality
sexuell	sexual
sexuella	sexual
sexuellt	sexual
sfären	sphere
shahen	shah
shakespeare	shakespeare
shakespeares	shakespeare
sharia	sharia
sheen	sheen
sibirien	siberia
sicilien	sicily
sida	page
sidan	page
side	side
sidor	pages
sidorna	the pages
sierra	sierra
siffra	figure
siffran	figure
siffror	figures
siffrorna	figures
sig	to
sigmund	sigmund
signaler	signals
signifikant	significant
sikt	term
silver	silver
simmons	simmons
simning	swimming
simon	simon
simpson	simpson
simpsons	simpsons
sin	its
sina	their
sinatra	sinatra
singapore	singapore
singapores	singapore
singel	single
singeln	single
singer	singer
singlar	singles
singlarna	singles
sinne	mind
sir	sir
sist	last
sista	last
siste	last
sistnämnda	last
site	site
sitt	his
sitta	sit
sittande	sitting
sitter	serve
situation	situation
situationen	situation
situationer	situations
siv	siv
sixx	sixx
sju	seven
sjuk	ill
sjuka	disease
sjukdom	disease
sjukdomar	diseases
sjukhus	hospital
sjukhuset	hospital
sjukvård	healthcare
sjunde	seventh
sjunga	sing
sjunger	sings
sjunka	decrease
sjunkande	sinking; decreasing
sjunker	flag
sjunkit	sunk
själ	soul
själen	soul
själv	self
själva	self
självbiografi	autobiography
självklart	course
självmord	suicide
självstyrande	autonomous
självstyre	autonomy
självständig	independent
självständiga	independent
självständighet	autonomy
självständigheten	independence
självständigt	independent
självt	itself
sjätte	sixth
sjö	lake
sjöar	lakes
sjöarna	lakes
sjöfart	shipping
sjöfarten	shipping
sjögren	sjögren
sjön	lake
sjöng	sang
sjönk	decreased
sjöss	sea
sk	so called
ska	should
skabb	scabies
skada	damage
skadad	damaged
skadade	damaged
skadades	wounded
skadan	damage
skadas	damaged
skadliga	deleterious
skador	damage
skadorna	damage
skaffa	get
skaffade	provided
skal	shell
skala	scale
skalan	scale
skalet	shell
skall	shall
skalv	quake
skalvet	quake
skandinavien	scandinavia
skandinaviska	scandinavian
skapa	create
skapad	created
skapade	created
skapades	created
skapande	creative
skapandet	creation
skapar	creates
skapare	creator
skapas	creates
skapat	designed
skapats	created
skapelse	creation
skara	city in south-central sweden (uppland)
skarp	sharp
skarsgård	skarsgård
skatt	tax
skatter	taxes
ske	happen
skedde	was
skede	phase
skelett	skeleton
skepp	ship
skeppen	the ships
skeppet	ship
sker	done
skett	occurred
skick	condition
skicka	send
skickade	sent
skickades	sent
skickar	sends
skickas	sent
skicklig	skillful
skiftande	changing
skikt	layer
skilda	different
skilde	divided
skildes	separated
skildrar	describes
skildras	is depicted
skildringar	description
skilja	distinguish
skiljas	separated
skiljer	different
skiljs	separated
skillnad	difference
skillnaden	difference
skillnader	differences
skillnaderna	differences
skilsmässa	divorce
skiva	disc
skivan	disc
skivbolag	label
skivbolaget	label
skivkontrakt	record deal
skivor	plates
skivorna	the records
skjuta	delay
skjuten	shot
skjuter	shoots
skog	forest
skogar	forests
skogarna	forests
skogen	woods
skola	school
skolan	school
skolgång	schooling
skolor	schools
skolorna	schools
skor	shoes
skorpan	crust
skotsk	scottish
skotska	scottish
skott	shot
skottland	scotland
skov	relapse
skrev	wrote
skrevs	august
skrift	writing
skriften	no.
skrifter	writings
skrifterna	scriptures
skriftliga	written
skriva	write
skrivas	printed
skriven	written
skriver	write
skrivet	written
skrivit	written
skrivits	written
skrivna	written
skrivs	printed
skräck	horror
skuggan	the shadow
skuld	debt
skulden	debt
skulder	liabilities
skull	sake
skulle	would
skulptur	sculpture
sky	sky
skydd	protection
skydda	protect
skyddade	protected
skyddar	protection
skyddas	protected
skyldig	guilty
skyskrapor	high rise buildings; sky scrapers
skäl	reason
skär	will
skära	cut
skärgård	archipelago
skådespelare	actor
skådespelaren	actor
skådespelarna	actors
skådespelerska	actress
skåne	skåne
skånes	scania's
skånska	skånska
skönhet	beauty
skönlitteratur	fiction
sköt	shot
sköta	handle
sköter	handles
sköts	shot
sköttes	operated
slag	kind
slaget	stroke
slagit	beaten
slags	kind
slavar	slaves
slaveriet	slavery
slaviska	slavic
slidan	vaginal
slipknot	slipknot
slippa	avoid
slog	beat
slogs	fought
slott	castle
slottet	castle
slovakien	slovakia
slovenien	slovenia
slovenska	slovenian
slut	final
sluta	stop
slutade	finished
slutar	ends
slutat	longer
slutet	end
slutgiltiga	final
slutliga	final
slutligen	at last
slutsats	conclusion
slutsatsen	the conclusion
slutsatser	conclusions
släkt	family
släkten	the family
släktet	genus
släkting	relative
släktingar	relatives
släktskap	relationship
släppa	drop
släppas	released
släpper	release
släpps	released
släppt	released
släppte	released
släpptes	released
släppts	released
slå	beat
slår	beat
slås	switched
slåss	fight
slöt	closed
slöts	concluded
sm	s-m
smak	taste
smaken	flavor
smala	narrow
smallwood	smallwood
smeknamn	nickname
smeknamnet	nickname
smguld	swedish championship gold
smith	smith
smitta	infection
smycken	jewlery
smält	melted
smärta	pain
små	small
småland	smaland
smålands	smaland's
småningom	gradually
snabb	fast
snabba	rapid
snabbare	faster
snabbast	fastest
snabbaste	fastest
snabbt	quickly
snarare	rather
snarast	rather
snart	soon
snitt	cut
snittet	section
snus	snuff
snuset	snuff
snö	snow
social	social
sociala	social
socialdemokrater	social
socialdemokraterna	members of the social democracy
socialdemokratiska	socialist
socialism	socialism
socialismen	socialism
socialister	socialists
socialistisk	socialist
socialistiska	socialist
socialistiskt	socialist
socialt	social
socken	parish
socker	sugar
sofia	sofia
sofie	sofie
sokrates	socrates
sol	sun
soldat	soldier
soldater	troops
soldaterna	soldiers
solen	sun
solens	the sun
solljus	sunlight
soloalbum	solo album
solsystem	solar system
solsystemet	solar system
solsystemets	solar system
solvinden	the solar wind
som	as
somalia	somalia
somliga	some
sommar	summer
sommaren	summer
sommarspelen	summer games
sommartid	summer-time
somrar	summers
somrarna	summers
son	son
sonen	son
sony	sony
sorg	grief
sorter	varieties
sorters	kinds
sorts	variety
soul	soul
sound	sound
soundtrack	soundtrack
south	south
sover	sleep
sovjet	soviet
sovjetisk	soviet
sovjetiska	soviet
sovjetunionen	soviet union
sovjetunionens	soviet union
spaniel	spaniel
spanien	spain
spaniens	spain
spanjorerna	the spaniards
spannmål	cereals
spansk	spanish
spanska	spanish
sparken	park
sparta	sparta
spears	spears
special	compare
specialiserade	specialized
speciell	special
speciella	special
specifik	specific
specifika	specific
specifikt	specifically
speglar	mirrors
spektrum	spectrum
spektrumet	spectrum
spekulationer	speculations
spel	game
spela	play
spelad	played
spelade	played
spelades	filmed
spelar	play
spelare	player
spelaren	player
spelarna	players
spelas	played
spelat	played
spelats	recorded
spelen	games
spelet	game
spelfilmer	movies
spelning	gig
spelningar	shows
spelningen	show
spets	edge; top
spetsen	edge; top
spetshundar	tip of dogs
spindlar	spiders
spindlingar	cortinarius
splittrades	split
spontant	spontaneously
sport	sports
sporten	port
sporter	sports
spotify	spotify
spred	spread
spreds	spread
sprida	spread
spridas	disseminated
spridd	scattered
spridda	spread
sprider	spreading
spridit	spread
spridning	diffusion
spridningen	spreading
sprids	spreads
springer	runs
springsteen	springsteen
springsteens	springsteens
sprit	liqeur
spritt	spread
språk	language
språkbruk	parlance
språken	languages
språket	language
språkets	language
språkliga	linguistic
spänner	range
spänning	voltage
spänningar	tensions
spänningen	voltage
spår	track
spåra	track
spåras	trace
spåren	the tracks
spårvagnar	trams
sr	sr
sri	sri
ss	ss
st	saint
stabil	stable
stabila	stable
stabilitet	stability
stad	city
staden	city
stadens	city
stadigt	stable
stadion	stadium
stadium	stage
stadsbild	cityscape
stadsdel	district
stadsdelar	districts
stadsdelarna	districts
stadsdelen	neighborhood
stadshus	town hall
stadskärna	center
stadskärnan	center
stadsparken	city park
staffan	staffan
stalin	stalin
stalins	stalin
stallone	stallone
stam	tribe
stammar	tribes
stammarna	tribes
stan	town
stand	stand
standard	standard
stanley	stanley
stanna	stay
stannade	stayed
stannar	stop
stark	strong
starka	strong
starkare	stronger
starkast	strongest
starkaste	strongest
starkt	strong
start	start
starta	start
startade	started
startades	started
startar	start
startat	started
starten	start
stat	state
state	state
statens	state
stater	states
staterna	states
staternas	states
states	states
station	station
stationen	station
stationer	stations
statistik	statistics
statistiska	statistical
statlig	state
statliga	governmental
statligt	state
stats	state
statschef	head of state
statschefen	head of state
statskupp	coup
statsmakten	the government
statsminister	prime minister
statsministern	prime minister
statsreligion	state religion
statsskick	government
statsöverhuvud	head of state
status	status
staty	statue
statyn	statue
stavning	spelling
stavningen	spelling
stefan	stefan
steg	step
steget	step
sten	stone
stenar	stones
stephen	stephen
steve	steve
steven	steven
stewart	stewart
stieg	stieg
stift	pin
stiftelsen	foundation
stig	stig
stiga	rise
stigande	rising
stiger	rising
stilar	styles
stilen	style
stilla	still
stimulans	stimulation
stimulera	stimulate
stimulerar	stimulates
stjäla	steal
stjärna	star
stjärnan	star
stjärnans	star
stjärnor	stars
stjärnornas	the star's
stockholm	stockholm
stockholms	stockholm's
stod	was
stoft	dust
stol	chair
stolpiller	suppository
stommen	body
stop	stop
stopp	stop
stoppa	stop
stoppade	stop
stor	big
stora	large
storbritannien	uk
storbritanniens	uk
store	great
stores	the great
storhetstid	greatness
storkors	the grand cross
storlek	size
storleken	size
storm	storm
stormakt	great power
stormakter	powers
stormakterna	great powers
stormaktstiden	great power
storstäder	metropolises
stort	large
stortorget	stortorget
story	story
straff	penalty
straffet	penalty
strand	beach
stranden	beach
strategiska	strategic
stratton	stratton
strax	just
streck	line
stred	fought
street	street
stress	stress
stressorer	stressors
strid	fight
strida	conflict
stridande	fighting
striden	fight
strider	battles
striderna	battles
stridigheter	oppositions
strikt	strict
strikta	strict
strindberg	strindberg
strindbergs	strindberg's
struktur	structure
strukturen	structure
strukturer	structures
sträckan	the distance
sträcker	extend
sträckor	routes
sträckte	extended
stränder	beaches
sträng	string
stränga	severe
strävan	endeavor
strävar	strives
strävhårig	hispid
strålning	radiation
strålningen	radiation
ström	current
strömmar	flow
strömmen	current
strömning	flow
strömningar	sentiments
stuart	stuart
student	student
studenter	students
studenterna	students
studera	study
studerade	studied
studerar	study
studeras	studied
studerat	studied
studie	study
studien	study
studier	studies
studierna	studies
studiet	study
studio	studio
studioalbum	studio album
studioalbumet	studio album
studion	studio
studios	studios
stulna	stolen
stund	while
stundom	sometimes
stupade	fallen
sture	sture
stycke	piece
stycken	pieces
styr	control
styra	steer
styrande	rulers
styras	controlled
styrde	ruled
styrdes	controlled
styre	rule
styrelse	board
styrelsen	board of directors
styrelseskick	government
styret	gate
styrka	strength
styrkan	strength
styrkor	strenghts
styrkorna	forces
styrs	controlled
städer	cities
städerna	urban
ställa	put
ställas	prepared
ställde	set
ställdes	prepared
ställe	place
ställen	spots; places
ställer	down
stället	instead
ställning	position
ställningar	positions
ställningen	score
ställs	is
ställt	set
stämma	meeting
stämmer	correct
ständerna	the cities
ständig	permanent
ständiga	standing
ständigt	constant
stänga	close
stängdes	closed
stängt	closed
stärka	strengthen
stärkelse	starch
stärkte	strengthened
stärktes	strengthened
stätta	stile
stå	stand
stående	standing
stål	steel
stålgemenskapen	steel community
stånd	stand
ståndpunkt	position
står	standing
stått	stood
stöd	support
stödde	supported
stöder	supports
stödet	aid
stödja	support
stödjer	supports
stöds	supported
störningar	disorders
större	major
störst	most
största	largest
störta	rush
störtades	overthrew
stöter	run
stött	supported
stövare	beagle
substantiv	noun
successivt	successively
succé	success
sudan	sudan
sugga	sow
sultanen	sultan
summa	amount
summan	sum
summer	sommar
sun	sun
sund	sound
sundsvall	sundsvall
sundsvalls	sundsvall
super	super
supportrar	supporters
sur	sour
susan	susan
sushi	sushi
sutra	sutra
suttit	sat
suverän	sovereign
suveräna	sovereign
suveränitet	sovereignty
sv	south west
svag	weak
svaga	weak
svagare	weaker
svagt	low
svar	response
svarade	accounted (for); answered
svarar	responds
svart	black
svarta	black
svartån	svartån
svavel	sulphur
svealand	svealand
sven	sven
svensk	swedish
svenska	swedish
svenskan	swedish
svenskans	swedish language
svenskar	swedish
svenskarna	swedish
svenske	swedish
svenskspråkiga	swedish speaking
svenskt	swedish
svensson	smith
sverige	sweden
sverigedemokraterna	sweden democrats
sveriges	sweden
svt	svt
svält	starvation
svärd	sword
svår	difficult
svåra	difficult
svårare	difficult
svårigheter	difficulties
svårt	difficult
swahili	swahili
swan	swan
sweden	sweden
swedish	swedish
sweet	söt
swift	swift
syd	south
sydafrika	south africa
sydafrikanska	south african
sydafrikas	south africa
sydamerika	south america
sydeuropa	southern europe
sydkorea	south korea
sydliga	southern
sydligaste	southernmost
sydost	south east
sydostasien	south east asia
sydstaterna	the southern states
sydväst	southwest
sydvästra	southwest
sydöst	south east
sydöstra	south east
syfta	aim
syftade	alluded to
syftar	refers
syfte	purpose
syften	purpose
syftet	purpose
symbol	symbol
symbolen	symbol
symboler	symbols
symboliserar	symbolizes
symbolisk	symbolic
symptom	symptom
symptomen	symptoms
symtom	symptoms
symtomen	symptoms
syn	sight
synd	sin
synder	sins
syndrom	syndrome
synen	sight
synes	seems to
synliga	visible
synligt	visible
synnerhet	especially
synnerligen	remarkably; particularly
synonymt	synonymously
syns	visible
synsätt	approach
synsättet	approach
syntes	showed
synvinkel	angle
syre	oxygen
syret	oxygen
syrgas	oxygen
syrien	syria
syskon	siblings
sysselsätter	employs
system	system
systematik	systematic
systematiska	systematic
systematiskt	systematic
systemet	system
systems	systems
syster	sister
systrar	sisters
säga	say
sägas	said
säger	says
sägs	how
säker	items
säkerhet	security
säkerheten	safety
säkerhetspolitik	security
säkerhetsråd	security
säkerhetsrådet	security
säkert	securely
säkra	secure
sälja	sell
säljande	selling
säljas	sold
säljer	selling
säljs	sold
sällan	rare
sällskap	company
sällskapet	society
sällskapshundar	pet dogs
sällsynt	rare
sällsynta	rare
sämre	poor
sämsta	worst
sända	send
sändas	broadcast
sände	sent
sändebud	messenger
sänder	sends
sändes	sent
sänds	sends
sänka	lower
sänker	lower
sänktes	reduced
särdrag	feature
särskild	special
särskilda	specific
särskilt	particulary
säsong	season
säsongen	season
säsongens	season
säsonger	seasons
säsongerna	seasons
säte	seat
sätt	way
sätta	put
sättas	added
sätter	puts
sättet	way
sätts	added
så	so
sådan	such
sådana	such
sådant	such
såg	saw
sågs	observed
sålda	sold
sålde	sold
såldes	was
således	thus
sålt	sold
sålts	sold
sålunda	thus
sång	singing
sångare	singer
sångaren	singer
sången	the song
sånger	songs
sångerna	songs
sångerska	singer
sår	wound
såsom	as
såväl	both
söder	south
söderut	south
södra	southern
söka	search
söker	searching
sökt	searched
sökte	searched
sömn	sleep
söndagen	sunday
sönder	broken
söner	sons
t	t
ta	take
tabell	chart
tabellen	table
tacitus	tacitus
tack	thanks
tackade	accepted
tag	while
tagen	taken
taget	time
taggar	spikes
tagit	taken
tagits	taken
taiwan	taiwan
taket	the roof
takt	rate
taktik	tactics
tala	speak
talade	spoke
talades	spoken
talang	talent
talanger	talents
talar	speaks
talare	speaker
talas	spoken
talat	spoken
talen	numbers
talet	the number
talets	century
talman	president
talmannen	president
talrika	numerous
tankar	thoughts
tanke	thought
tanken	thought
tanzania	tanzania
tappade	lost
tappar	drop
tar	takes
tas	is
taube	taube
taubes	taubes
taylor	taylor
te	tea
team	team
teater	theater
teatern	theater
teatrar	theaters
tecken	sign
tecknade	signed
tecknet	sign
ted	ted
teddy	teddy
tegel	brick
teknik	technique
tekniken	art
tekniker	technician
teknisk	technical
tekniska	technology
tekniskt	technical
teknologi	technology
telefon	phone
telefonen	phone
telegram	telegram
television	television
tema	theme
teman	themes
tempel	temple
temperatur	temperature
temperaturen	temperature
temperaturer	temperature
tempererat	temperature
templet	temple
tendens	tendency
tendenser	tendencies
tenderar	tend
tenn	tin
tennessee	tennessee
tennis	tennis
tennisspelare	tennis
teologi	theology
teologiska	theological
teoretiker	theorists
teoretisk	theoretical
teoretiska	theoretical
teoretiskt	theoretical
teori	theory
teorier	theories
teorin	theory
termen	term
termer	terms
terminologi	terminology
terrier	terrier
territoriella	territorial
territorier	territories
territorierna	territories
territoriet	territory
territorium	territory
terror	terror
terrorism	terrorism
terrorismen	terrorism
terrorister	terrorists
terry	terry
terräng	terrain
tesla	tesla
teslas	tesla's
test	test
testamente	testament
testamentet	testament
tex	for example
texas	texas
text	text
texten	text
texter	texts
texterna	texts
th	th
thailand	thailand
than	than
that	that
thc	thc
the	the
theodor	theodor
theta	theta
they	they
thierry	thierry
thomas	thomas
thriller	thriller
thåström	thåström
tibet	tibet
tid	time
tiden	time
tidens	time's
tider	times
tiderna	times
tiders	times
tidig	early
tidiga	early
tidigare	earlier
tidigast	the earliest
tidigt	early
tidning	newspaper
tidningar	magazines
tidningarna	papers
tidningen	newspaper
tidpunkt	time
tidpunkten	time
tids	time
tidskrift	journal
tidskriften	journal
tidskrifter	periodicals
tidszon	zone
tidszoner	time zones
tidvis	times
tiger	tiger
tigern	tiger
tigrar	tigers
till	to
tillbaka	back
tillbehör	accessory
tillbringade	spent
tillbringar	spends
tilldelades	awarded
tilldelas	awarded
tilldelats	assigned
tillfälle	occasion
tillfällen	occasion
tillfället	currently
tillfällig	temporary
tillfälliga	temporary
tillfälligt	temporarily
tillgänglig	available
tillgängliga	available
tillgängligt	available
tillgång	access
tillgångar	assets
tillgången	access
tillhandahåller	provides
tillhör	belonging to
tillhöra	belong
tillhörande	associated
tillhörde	belonged
tillhörighet	belonging
tillhört	belonged
tillika	also
tillkom	advent
tillkommer	will
tillkommit	accured
tillkomst	advent
tillkännagav	announced
tillräcklig	enough
tillräckliga	sufficient
tillräckligt	enough
tills	until
tillsammans	together
tillstånd	state
tillståndet	state
tillsätts	added
tilltagande	increasing
tillträdde	took
tillträde	access
tillvaron	existence
tillverka	manufacture
tillverkade	manufactured
tillverkar	makes
tillverkare	manufacturer
tillverkas	manufactured
tillverkning	production
tillverkningen	production
tillväxt	growth
tillväxten	growth
tilly	tilly
tillägg	addition
tillämpa	applying
tillämpar	applying
tillämpas	applied
tillämpningar	applications
tillät	allowed
tilläts	allowed
tillåta	allow
tillåtelse	permission
tillåter	allow
tillåtet	allowed
tillåtna	allowed
tillåts	allowed
tim	h
time	time
timmar	hours
timme	hour
tina	thaw
ting	things
tingslag	leet
tintin	tintin
tio	ten
tionde	tenth
tiotusentals	tens of thousands
titanic	titanic
titanics	titanic
titel	title
titeln	title
titlar	titles
titta	watch
tittar	looking; viewing; viewer
tittarna	viewers
tjeckien	czech
tjeckiska	czech
tjeckoslovakien	czechoslovakia
tjugo	twenty
tjäna	serve
tjänade	earned
tjänar	earns
tjänare	servant
tjänst	service
tjänstemän	officials
tjänsten	service
tjänster	services
tobak	tobacco
tobias	tobias
tog	took
togs	was
tokyo	tokyo
tolerans	tolerance
tolfte	twelth
tolka	interpret
tolkade	interpreting
tolkar	interprets
tolkas	interpreted
tolkats	interpreted
tolkien	tolkien
tolkiens	tolkien
tolkning	interpretation
tolkningar	interpretations
tolkningen	interpretation
tolv	twelve
tom	empty
tomas	tomas
tomma	empty
tomt	empty
ton	t
tongivande	influential
tony	tony
top	top
topp	top
toppade	topped
toppar	tops
toppen	top
tor	thu
torah	torah
torbjörn	torbjorn
torde	should
torg	square
torget	square
torka	dry
torn	tower
tornen	towers
tornet	tower
toronto	toronto
torra	dry
torres	torres
torrt	dry
torsten	torsten
tortyr	torture
tosh	tosh
total	total
totala	total
totalt	total
tottenham	tottenham
tour	tour
toy	toy
tradition	tradition
traditionell	traditional
traditionella	traditional
traditionellt	traditional
traditionen	the tradition
traditioner	traditions
traditionerna	traditions
trafik	traffic
trafiken	traffic
trafikerade	trafficked
trafikerar	traffic
trafikeras	trafficked
trakten	area
transeuropeiska	ten
transkription	transcript
transport	transport
transporter	transport
transportera	transport
transporterar	carrying
transporteras	transported
tre	three
tredje	third
tredjedel	third
tredjedelar	thirds
tree	tree
treenigheten	trinity
treenighetsläran	the trinity
trend	trend
trenden	trend
trettio	thirty
trettioåriga	13 year olds
tretton	thirteen
trey	trey
triangel	triangle
triangeln	triangle
triangelns	triangle
trianglar	traingles
trigonometriska	trigonometric
trinidad	trinidad
tro	believe
trodde	thought
troende	faithful
troligen	probably
troligt	likely
troligtvis	probably
tron	faith
tronen	the throne
tronföljare	heir
tropisk	tropical
tropiska	tropical
tropiskt	tropical
tror	think
tros	belived
trosbekännelsen	creed
trossamfund	religious community
trots	although
trotskij	trotskij
truman	truman
trummis	drummer
trummisen	drummer
trummor	drums
trupp	troops
trupper	troops
trupperna	troops
tryck	print
trycket	pressure
tryckta	printed
trycktes	printed
trä	wood
träd	tree
träda	fallow
trädde	entry
träffa	hit
träffade	met
träffades	met
träffar	results
träffas	meet
träffat	met
tränade	trained
tränare	coach
tränaren	coach
tränga	push (aside)
tränger	forces forward
träning	exercise
trådlös	wireless
trött	tired
tsar	tsar
tsaren	czar
tsunami	tsunami
tsunamier	tsunamis
tum	inch
tung	heavy
tunga	tongue
tungt	heavy
tunisien	tunisia
tunn	thin
tunna	thin
tunnel	tunnel
tunnelbana	subway
tunnelbanan	subway
tunnlar	tunnels
tupac	tupac
tur	lucky
turism	tourism
turismen	tourism
turister	tourists
turistmål	tourist destination
turkar	turks
turkarna	turks
turkiet	turkey
turkiets	turkey
turkisk	turkish
turkiska	turkish
turner	tournament
turnera	tour
turnerade	toured
turneringen	tournament
turné	tour
turnéer	tours
turnén	tour
tusen	thousands
tusentals	thousands
tv	tv
tvfilm	tv-movie
tvinga	force
tvingade	forced
tvingades	forced
tvingas	forced
tvingats	forced
tvister	disputes
tvkanaler	tv channels
tvprogram	tv program
tvserie	tv series
tvserien	tv series
tvserier	tv series
tvskådespelare	tv actor
tvungen	forced
tvungna	had
tvärtom	on the contrary
två	two
tvåa	second
twilight	twilight
ty	for
tycker	think
tyckte	thought
tycktes	seemed
tyder	indicates
tydlig	clear
tydliga	clear
tydligt	clear
tyngre	heavier
typ	type
typen	type
typer	types
typerna	types
typisk	typical
typiska	typical
typiskt	typical
tysk	german
tyska	german
tyskar	germans
tyskarna	germans
tyske	german
tyskland	germany
tysklands	germany
tyskt	german
tyst	silent
tyvärr	unfortunately
täcka	cover
täcker	covers
täcks	covered
täckt	covered
tämligen	rather
tänder	teeth
tänderna	teeth
tänka	think
tänkande	thinking
tänkandet	thinking
tänkare	thinker
tänker	thinking
tänkt	thought
tänkte	thought
tät	close
täta	close
tätbefolkade	densely populated
tätort	urban
tätorten	conurbation
tätorter	urban
tätt	tight
tävla	compete
tävlade	competed
tävling	contest
tävlingar	competitions
tävlingen	competition
tåg	train
tågen	trains
tåget	train
tål	stand
u+	u +
udda	odd
uefa	uefa
uefacupen	the uefa champions league
uganda	uganda
ugandas	uganda
uggla	owl
ugglas	ugglas
uk	uk
ukraina	ukraine
ukrainas	ukraine
ukrainska	ukrainian
ulf	ulf
ullevi	ullevi
ulrich	ulrich
ultraviolett	ultraviolet
umgänge	intercourse
und	und
undan	away
undantag	exception
undantaget	except
under	during
underart	subspecies
underarten	subspecies
underarter	subspecies
undergång	doom
underhåll	support
underhållning	entertainment
underjordiska	underground
underliggande	underlying
underlätta	facilitate
underlättar	make it easier
underordnade	subordinates
undersöka	study
undersökning	investigation
undersökningar	studies
undersökte	examined
undertecknades	signed
underverk	wonder
undervisade	taught
undervisning	teaching
undervisningen	teaching
undre	lower
undvika	avoid
undviker	avoid
unesco	unesco
unescos	unesco
ung	young
unga	young
ungar	kids
ungarna	kids
ungdom	youth
ungdomar	adolescents
unge	young
ungefär	approximately
ungern	hungary
ungerns	hungary
ungerska	hungarian
uniform	uniform
unik	unique
unika	unique
unikt	unique
union	union
unionen	union
unionens	union
universitet	university
universiteten	universities
universitetet	university
universum	universe
universums	universe
uno	uno
up	up
upp	up
uppbyggd	structured
uppbyggnad	construction
uppbyggt	structured
uppdelad	divided
uppdelade	broken
uppdelat	divided
uppdelning	division
uppdelningen	division
uppdrag	mission
uppdraget	assignment
uppe	up
uppehåll	rain
uppemot	up
uppenbarelse	revelation
uppenbarelser	revelations
uppfann	invented
uppfanns	invented
uppfatta	perceive
uppfattade	perceived
uppfattar	perceive
uppfattas	perceived
uppfattning	understanding
uppfattningar	perceptions
uppfattningen	view
uppfinnare	inventor
uppfinningar	inventions
uppfostran	upbringing
uppfylla	meet
uppfyller	fulfills
uppföljare	sequel
uppförande	conduct
uppfördes	was constructed
uppgav	stated
uppger	state
uppges	reported
uppgick	total
uppgift	task
uppgiften	task
uppgifter	tasks
uppgifterna	information
uppgörelse	settlement
upphov	rise
upphovsman	author
upphovsrätt	copyright
upphovsrätten	copyright
upphörde	ceased
upphört	ceased
uppkallad	named
uppkom	arose
uppkommer	occur
uppkommit	arisen
uppkomst	origin
uppkomsten	appearance
upplaga	edition
upplagan	the edition
upplagor	editions
uppleva	experience
upplevde	experiences
upplevelse	experience
upplevelser	experiences
upplever	experience
upplysning	information
upplysningen	the enlightenment
upplysningstiden	enlightenment
upplösning	resolution
upplösningen	disbandment
upplöstes	dissolved
uppmanade	called
uppmaning	call
uppmuntrade	encouraged
uppmärksamhet	attention
uppmärksammad	noticed
uppmärksammade	attention
uppmärksammades	attention
uppmärksammat	attention
uppnå	achieve
uppnådde	achieved
uppnår	achieve
uppnås	obtained
uppnått	met
upprepade	repeated
uppror	rebellion
upproret	uprising
upprustning	renovation
upprätta	establish
upprättade	prepared
upprättades	established
upprättandet	establishment
upprättas	established
upprätthålla	maintain
upprätthåller	maintains
uppsala	uppsala
uppskatta	appreciate
uppskattad	appreciated
uppskattade	estimated
uppskattades	estimated
uppskattar	estimates
uppskattas	estimated
uppskattning	appreciation
uppskattningar	estimates
uppskattningsvis	estimated
uppslagsordet	entry word
uppslagsverk	encyclopedia
uppstod	arose
uppstå	develop
uppståndelse	resurrection
uppstår	occur
uppstått	occurred
uppsving	boost
uppsättning	set
upptagen	occupied
upptar	occupies
uppträda	act
uppträdande	performance
uppträdde	occurred
uppträder	occur
upptäcka	discover
upptäcker	discoveries
upptäcks	detected
upptäckt	discovered
upptäckte	discovered
upptäckten	discovery
upptäckter	discoveries
upptäcktes	detected
uppvisade	showed
uppvisar	shows
uppvärmning	heating
uppvärmningen	heating
uppväxt	childhood
uppåt	up
ur	from
uralbergen	the ural mountains
uran	uranium
urin	urine
urskilja	distinguish
ursprung	origin
ursprunget	origin
ursprungliga	original
ursprungligen	originally
ursprungsbefolkning	native population
ursprungsbefolkningen	the native population
ursäkt	excuse
uruguay	uruguay
urval	selection
usa	usa
usama	usama
usas	usa
ut	out
utan	without
utanför	outside
utbildad	educated
utbildade	educated
utbildning	training
utbildningen	training
utbredd	widespread
utbredda	widespread
utbredning	spread
utbrett	spread
utbrott	outbreak
utbröt	erupted
utbud	range
utbyggda	expanded
utbyggnad	development
utbyggt	expanded
utbyte	exchange
utdelades	awarded
utdöda	extinct
ute	out
uteslutande	exclusively
utformade	formed
utformning	layout
utformningen	the layout
utfärdade	issued
utför	perform
utföra	perform
utföras	performed
utförd	performed
utförda	executed
utfördes	performed
utförs	performed
utfört	performed
utgavs	issued
utgick	started
utgifter	expenditure
utgiven	published
utgivna	issued
utgivningen	release
utgjorde	was
utgjordes	make up
utgångspunkt	starting point
utgår	deleted
utgåva	edition
utgåvan	edition
utgåvor	editions
utgör	constitutes
utgöra	represent
utgörs	consists of
utifrån	from
utkanten	edge
utkom	published
utkämpades	fought
utlandet	abroad
utlopp	outlet
utländsk	foreign
utländska	foreign
utlänningar	foreigners
utlösa	trigger
utlösning	release
utlöste	triggered
utmed	along
utmärkande	characteristic
utmärkelsen	award
utmärkelser	awards
utmärker	characterizes
utmärks	characterized
utmärkt	excellently
utnyttja	use
utnyttjade	utilized
utnyttjar	using
utnyttjas	utilized
utnämndes	named
utom	except
utomeuropeiska	non-european
utomlands	abroad
utomliggande	external; ex-territorial
utomstående	outsider
utredning	investigation
utredningen	investigation
utrikes	foreign
utrikesminister	minister of foreign affairs
utrikespolitik	foreign policy
utrikespolitiken	foreign policy
utrikespolitiska	foreign policy
utropade	exclaimed
utropades	proclaimed
utrotning	extinction
utrustning	equipment
utrymme	space
utsatt	exposed
utsatta	exposed
utsattes	subjected
utse	appoint
utsedd	designated
utseende	appearance
utser	appoints
utses	designated
utskott	committee
utsläpp	emissions
utspelar	set
utsträckning	extent
utställning	exhibition
utsätts	exposed
utsåg	appointed
utsågs	was
utsöndras	secrete
uttal	pronunciation
uttalade	pronounced
uttalande	statement
uttalanden	statements
uttalas	pronounced
uttalat	pronounced
uttalet	the pronounciation
uttryck	expression
uttrycka	express
uttrycker	express
uttrycket	the expression
uttryckligen	explicitly
uttryckt	expressed
uttryckte	expressed
utvalda	selected
utveckla	develop
utvecklad	developed
utvecklade	developed
utvecklades	developed
utvecklandet	development
utvecklar	develops
utvecklas	develop
utvecklat	developed
utvecklats	developed
utveckling	development
utvecklingen	development
utvidgade	expanded
utvidgning	enlargement; expansion
utvinna	extract
utvinns	extracted
utvisning	penalty
utåt	outwardly
utökade	extended
utökat	expanded
utöva	exercise
utövade	exercised
utövar	exercise
utövas	is practised
vacker	beautiful
vackra	beautiful
vad	what
vaginalt	vaginal
vagn	wagon
vagnar	wagons
val	choice
valborg	valborg
vald	selected
valda	selected
valde	crowned
valdes	elected
valen	elections
valet	election
valla	wax
valley	valley
vallhund	herder
valrörelsen	election
valt	selected
valuta	currency
valutan	currency
vampyr	vampire
vampyren	vampire
vampyrer	vampire
van	van
vana	familiar
vandrar	wanders
vanföreställningar	delusions
vanlig	common
vanliga	usual
vanligare	common
vanligast	common
vanligaste	most common
vanligen	usually
vanligt	usual
vanligtvis	usually
vann	won
vanns	won
vapen	arms
vapnen	weapons
vapnet	force
var	where
vara	be
varade	lasted
varandra	each other
varandras	each others
varar	lasts
varav	which
vardagen	everyday
vardagliga	everyday
vardagligt	everyday
vardera	each
vare	to
varefter	whereafter
varelse	creature
varelser	creatures
varför	why
varg	wolf
vargar	wolves
vargen	wolf
variant	variant
varianten	variant
varianter	variants
varianterna	variants
variation	diversity
variationer	variations
variera	vary
varierade	varied
varierande	varying
varierar	varies
varierat	varied
varifrån	where
varit	been
varje	each
varken	neither
varm	warm
varma	hot
varmare	warmer
varmblod	warmblood
varmed	whereby
varmt	hot
varna	varna
varnade	warned
varning	warning
varor	goods
varpå	whereupon
vars	whose
varsin	each
vart	where
varuhus	department store
varv	turn
varvid	in which
vasa	vasa
vasaloppet	vasaloppet
vasas	vasa
vatikanstaten	vatican
vatten	water
vattendrag	water
vattenkraft	water power
vattenånga	steam
vattnet	water
vattnets	water
vd	ceo
vecka	week
veckan	the week
veckor	weeks
veckorna	weeks
vegas	vegas
velat	liked
vem	who
venedig	venice
venezuela	venezuela
venus	venus
verde	verde
verk	work
verka	act
verkade	seemed
verkan	effect
verkar	seems
verkat	acted
verken	plants
verket	plant
verklig	real
verkliga	real
verkligen	really
verklighet	reality
verkligheten	real
verksam	active
verksamhet	operation
verksamheten	business
verksamheter	operations
verksamma	active
verkställande	executive
verktyg	tool
vers	verse
versaillesfreden	treaty of versailles
version	version
versionen	release
versioner	versions
vet	know
veta	know
vete	wheat
vetenskap	science
vetenskapen	science
vetenskaplig	scientific
vetenskapliga	scientific
vetenskapligt	scientifically
vetenskapsmän	scientists
veto	veto
vhs	vhs
vi	we
via	via
vice	vice
vicepresident	vice
victor	victor
victoria	victoria
victoriasjön	lake victoria
vid	at
vida	far
vidare	further
video	video
videon	video
vidsträckta	broad
vidta	take
vietnam	vietnam
vietnamesiska	vietnamese
vietnamkriget	vietnam war
vietnams	vietnam
viggo	viggo
vii	vii
vika	fold
viken	gulf
viking	viking
vikingar	vikings
vikingarna	the vikings
vikingatiden	the viking age
vikt	weight
vikten	weight
viktig	important
viktiga	important
viktigare	important
viktigaste	important
viktigt	important
viktor	viktor
vila	rest
vilar	rest
vilda	wild
vilhelm	vilhelm
vilja	will
viljan	will
vilka	which
vilkas	whose
vilken	which
vilket	which
vill	want
villa	villa
ville	wanted
villkor	terms
villkoren	conditions
villor	villas
vimmerby	vimmerby
vin	wine
vincent	vincent
vinci	vinci
vind	wind
vindar	winds
vinden	the wind
vindkraft	wind
vindkraftverk	wind turbine
vingar	wings
vinkel	angle
vinkeln	angle
vinklar	angles
vinna	win
vinnare	winner
vinnaren	winner
vinner	wins
vinst	profit
vinsten	gain
vinster	profit
vinter	winter
vintergatan	milky way
vinterkriget	the winter war
vintern	winter
vinterspelen	winter games
vintertid	winter-time
vintrar	winters
vintrarna	winters
virginia	virginia
virus	virus
viruset	virus
vis	way
visa	show
visade	showed
visades	showed
visar	shows
visas	is shown
visat	found
visats	demonstrated
visby	visby
visdom	wisdom
vision	vision
visor	songs
viss	certain
vissa	some
visserligen	certainly
visst	certainly
visste	did
vista	vista
vistas	live
vistelse	stay
vit	white
vita	white
vitryssland	belarus
vitt	white
vittne	witness
vittnen	witnesses
vladimir	vladimir
vm	world championship
voddler	voddler
vojvodina	vojvodina
vojvodskap	voivodeship
vol	v
voltaire	voltaire
volvo	volvo
volym	volume
von	von
vore	would
vrida	turn
vulkaner	volcanoes
vulkaniska	volcanic
vulkanutbrott	vulcano eruption
vunnit	won
vuxen	adult
vuxit	grown
vuxna	adult
väckt	brought
väckte	aroused
väder	weather
vädret	weather
väg	way
vägar	ways
vägarna	paths
vägen	way
väger	weighs
vägg	wall
vägnät	road network
vägnätet	road network
vägrade	refused
vägrar	refuses
väl	selecting
väldet	empire
väldiga	immense
väldigt	very
välfärd	welfare
välgörenhet	charity
välja	select
väljas	selected
väljer	select
väljs	selected
välkänd	well-known
välkända	known
välmående	prosperous
välstånd	prosperity
vän	friend
vända	turn
vände	turned
vänder	face
vännen	the friend
vänner	friends
vänskap	friendship
vänster	left
vänstern	western
vänsterpartiet	left
vänstra	left
vänt	waiting
vänta	wait
väntade	waited
väntan	waiting
väntar	waiting
väntas	expected
väntat	expected
väpnad	armed
väpnade	armed
värd	host
värde	value
värdefulla	valuable
värden	values
värderingar	values
värdet	value
värld	world
världen	world
världens	the world
världsarv	world
världsarvslista	world heritage
världsbanken	world bank
världsdel	continent
världshälsoorganisationen	world health organization
världskrigen	the world wars
världskriget	world war
världskrigets	world war
världsliga	secular
världsrekord	world record
världsturné	world tour
värme	thermal
värmestrålningen	heat radiation
värmland	wermlandia
värmlands	new
värnplikt	military service
värnpliktiga	conscripted
värre	worse
värsta	worst
värt	worth
värvade	referred
väsen	entity
väsentligt	substantially
väska	bag
väst	west
västbanken	the west bank
västberlin	west berlin
väster	west
västerbottens	västerbottens
västergötland	västergötland
västerländsk	western
västerländska	western
västerut	west
västerås	västerås
västeuropa	western europe
västindien	caribbean
västkusten	the west coast
västlig	western
västliga	western
västmakterna	western powers
västra	western
västsahara	western sahara
västtyskland	west germany
västvärlden	west
väte	hydrogen
vätet	hydrogen
vätska	liquid
växa	grow
växande	growing
växer	grow
växjö	växjö
växt	plant
växte	grew
växter	plants
växterna	plants
växthuseffekten	the greenhouse effect
växthusgaser	vaxthusgaser
våg	wave
vågade	dared
vågen	the wave
våglängder	wavelengths
vågor	waves
våld	violence
våldet	violence
våldsam	violent
våldsamma	violent
våningar	levels
vår	spring
våra	our
vård	care
våren	spring
vårt	our
w	w
wagner	wagner
wahlgren	wahlgren
wailers	wailers
wales	wales
wall	wall
wallace	wallace
wallander	wallander
wallenberg	wallenberg
wallenstein	wallenstein
walt	walt
walter	walter
want	want
war	war
warhol	warhol
warner	warner
warszawa	warsaw
washington	washington
waterloo	waterloo
watson	watson
way	way
wayne	wayne
we	we
webbkällor	websources
webbplats	website
webbplatsen	website
webbplatser	websites
weber	weber
welsh	welsh
wembley	wembley
werner	werner
west	west
what	what
who	who
wien	vienna
wikipedia	wikipedia
wikipedias	wikipedia
wild	wild
wilde	wilde
wilhelm	wilhelm
will	will
william	william
williams	williams
willy	willy
wilson	wilson
wind	wind
winnerbäck	winnerbäck
winston	winston
without	without
wittenberg	wittenberg
wolfgang	wolfgang
works	works
world	world
wright	wright
x	x
xi	xi
xii	xii
xiis	xii
xis	the eleventh's
yngre	younger
yngsta	youngest
yngste	youngest
york	york
yorks	york
you	you
youtube	youtube
yta	surface
ytan	surface
ytterligare	further
ytterst	very; extremely
yttersta	furthest
yttre	outer
z	z
zach	zach
zagreb	zagreb
zanzibar	zanzibar
zarathustra	zarathustra
zeeland	zeeland
zeppelin	zeppelin
zeus	zeus
zink	zinc
zirkon	zircon
zlatan	zlatan
zon	zone
zonen	zone
zoner	zones
zuckerberg	zuckerberg
 cm	cm
 kilometer	kilometer
 km	kilometers
 kmh	km/h
 km²	km²
 meter	meter
 miljoner	million
 mm	millimeter
 procent	percent
  km²	km²
 °c	celsius
£m	million pounds
×	x
à	river
äga	own
ägande	owning
ägare	owner
ägda	run
ägde	took
ägdes	owned
äger	own
ägg	egg
ägna	spend
ägnade	spent
ägnar	spend time
ägs	owned
ägt	taken
äkta	genuine
äktenskap	marriage
äktenskapet	marriage
äldre	older
äldsta	oldest
äldste	elders
älg	moose
älgar	moose
älgen	elk; moose
älska	love
älskade	loved
älskar	love
ämbetsmän	officers
ämne	subject
ämnen	substances
ämnena	substances
ämnet	substance
än	than
ända	end
ändamål	purpose
ände	end
änden	end
ändra	change
ändrade	changed
ändrades	changed
ändrar	change
ändras	changed
ändrat	changed
ändringar	edit
ändå	still
änglar	angels
ängssyra	sorrel
ännu	yet
är	is
ära	oar
ärftliga	genetic
ärkebiskop	archbishop
ärkebiskopen	archbishop
äta	eat
äter	eat
ätten	the dynasty
ättlingar	descendants
även	also
äventyr	adventure
å	on
åka	go
åke	åke
åker	go
åkte	went
åland	Åland
ålands	Åland island's
ålder	age
åländska	Åland swedish
ån	from
ångest	anxiety
år	year
åren	years
årens	years
året	year
årets	year
århundraden	centuries
århundradena	centuries
århundradet	century
årig	old
åriga	-year
åring	age
årlig	annual
årliga	annual
årligen	annually
års	years
årsdag	anniversary
årstiderna	seasons
årsåldern	adult
årtionde	decade
årtionden	decades
ås	ridge
åsikt	opinion
åsikten	view
åsikter	opinions
åskådare	spectators
åstadkomma	achieve
åt	at
åtal	prosecution
åtalades	was prosecuted
åter	again
återfanns	was rediscovered
återfinns	found
återförening	reunion
återgick	went
återigen	again
återkom	return
återkommande	recurring
återkommer	returning
återkomst	return
återställa	resett
återstående	remaining
återstår	remains
återta	regain
återvända	return
återvände	returning
återvänder	returns
återvänt	returning
åtgärder	actions
åtminstone	at least
åtskilda	separated
åtskilliga	several
åtta	eight
åttonde	the eighth
ö	island
öar	islands
öarna	islands
öde	fate
ödleblad	houttuynia cordata
öga	eye
ögat	eye
ögon	eyes
ögonen	eyes
öka	increase
ökad	increased
ökade	increased
ökande	increasing
ökar	increases
ökat	increased
öken	desert
ökenråttor	gerbils
öknen	desert
ökning	increase
ökningen	increase
öl	beer
öland	öland
ölet	beer
ön	island
öns	island
önskade	desired
önskan	wish
önskar	desired
önskemål	requests
öppen	open
öppet	open
öppna	open
öppnade	opened
öppnades	opened
öppnat	opened
örebro	Örebro
öresund	sound
öron	ears
öronen	ears
öst	east
östafrika	east africa
östasien	east asia
östberg	Östberg
östberlin	east berlin
östblocket	east block
öster	east
östergötland	Östergötland
österrike	austria
österrikes	austria
österrikeungern	oster kingdom hungary
österrikiska	austrian
östersjön	baltic
österut	east
östeuropa	eastern europe
östfronten	eastern front
östman	Östman
östra	eastern
östtimor	east timor
östtyska	east german
östtyskland	east germany
östtysklands	east german
över	over
överallt	everywhere
överbefälhavare	commander
överens	agreed
överenskommelse	agreement
överensstämmer	conform
överföra	transfer
överföras	transfer
överföring	transfer
överförs	is transferred
övergav	abandoned
övergick	passed
övergrepp	abuse
övergripande	overall
övergå	pass
övergång	transition
övergången	transition
övergår	surpasses
överhuvudtaget	on the whole
överhöghet	supremacy
överleva	survive
överlevande	survivor; survivors; surviving
överlevde	survived
överlever	survives
överlevnad	survival
överlevt	survived
överlägset	superior
övernaturliga	supernatural
överraskande	surprisingly
övers	transl
översatt	translated
översikt	overview
överst	top
översvämningar	floodings
översättas	translated
översättning	translation
översättningar	translations
översättningen	translation
översätts	translated
övertala	persuade
övertalade	persuaded
övertog	took
övertogs	was taken
övertyga	convince
övervikt	overweight
övervägande	predominant
övre	upper
övrig	other
övriga	others
övrigt	other
